-------------------------------------------------------------------------------------------------------------
--
--  AVR Pipelined CPU TEST BENCH
--
--  This file contains the testbench for the Pipelined ATMEL AVR CPU. The testvectors generated for this testbench
--  originate from an AVR Simulator in Microchip Studio. The testvectors run through each of the operations
--  explained in the top level AVR CPU file and thoroughly checks each operation for correctness. 
--  
--  For each testvector (1 clock cycle) the following order of operations is performed:
-- 		the testbench will first load in data to the Program Data Bus
--      the testbench then checks the Program Address Bus immediately after loading in the program data bus
--      the testbench next waits until the rising edge of the CLK at which it ensures that DataDB is driven to 'Z'
--      the testbench then waits until the falling edge of the clock and then (if reading) loads data in the Data Data Bus
--  			      it also checks the Data Address Bus here for correctness
-- 		the testbench then waits for 0.1 us after falling edge and then checks the Data Data Bus (if writing) as well as the 
--                    read and write signals generated by the CPU for correctness
--
--  ** In order to test for pipelining, the test vector are shifted by 3 additional clock cycles. I.e. the first outputs
--     appear 4 clocks after sending in the first instruction through ProgDB. This means there are a total of 3 instructions
--     in process for the pipelined CPU at any given time. 
--
--  
--
--  Revision History:
--     02 Feb 23  Hector Wilson     Initial revision
--     10 Feb 23  Hector Wilson     Completed testbench
--     23 Feb 24  Hector Wilson     Added comments & updated test vectors
--     24 Feb 26  Hector Wilson     Updated test vectors
--     24 Feb 27  Hector Wilson     Updated test vectors
--     24 Mar 02  Hector Wilson     Updated test vectors
--     24 Mar 07  Hector Wilson     Updated test vectors
--     24 Feb 11  Hector Wilson     Updated test vectors
--     24 Feb 15  Hector Wilson     Updated test vectors
--     19 Mar 23  Hector Wilson     Updated comments
--     24 Mar 23  Hector Wilson     Updated TB for pipelined CPU
--     30 Mar 23  Hector Wilson     Updated comments
--
-------------------------------------------------------------------------------------------------------------
library opcodes;
use opcodes.opcodes.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all;    -- for uniform & trunc functions
use ieee.numeric_std.all;  -- for to_unsigned function

entity AVR_CPU_tb is
end AVR_CPU_tb;

architecture Behavioral of AVR_CPU_tb is
    component AVR_CPU 
        port ( 
	        ProgDB  :  in     std_logic_vector(15 downto 0);   -- program memory data bus
	        Reset   :  in     std_logic;                       -- reset signal (active low)
	        INT0    :  in     std_logic;                       -- interrupt signal (active low)
	        INT1    :  in     std_logic;                       -- interrupt signal (active low)
	        clock   :  in     std_logic;                       -- system clock
	        ProgAB  :  out    std_logic_vector(15 downto 0);   -- program memory address bus
	        DataAB  :  out    std_logic_vector(15 downto 0);   -- data memory address bus
	        DataWr  :  out    std_logic;                       -- data memory write enable (active low)
	        DataRd  :  out    std_logic;                       -- data memory read enable (active low)
	        DataDB  :  inout  std_logic_vector(7 downto 0)     -- data memory data bus
        );
    end component;

    -- set up test vectors
    type testarray is array (0 to 2764) of std_logic_vector(15 downto 0);
    type testarray2 is array (0 to 2764) of std_logic_vector(7 downto 0);

    -- Input Program Data Bus Vector
    constant ProgDataTest : testarray := (
		X"E203", X"9300", X"1000", X"1000", X"EF0F",
		X"9300", X"1000", X"1000", X"E001", X"9300",
		X"1000", X"1000", X"E000", X"9300", X"1000",
		X"1000", X"E415", X"9310", X"1000", X"1000",
		X"9100", X"1000", X"1000", X"9300", X"0900",
		X"0900", X"EF10", X"9310", X"1000", X"1000",
		X"9100", X"1000", X"1000", X"9300", X"0900",
		X"0900", X"E111", X"9310", X"1000", X"1000",
		X"9100", X"1000", X"1000", X"9300", X"0900",
		X"0900", X"E010", X"9310", X"1000", X"1000",
		X"9100", X"1000", X"1000", X"9300", X"0900",
		X"0900", X"EC0D", X"2EF0", X"92F0", X"1000",
		X"1000", X"E900", X"2EF0", X"92F0", X"1000",
		X"1000", X"E103", X"2EF0", X"92F0", X"1000",
		X"1000", X"E000", X"2EF0", X"92F0", X"1000",
		X"1000", X"EAAA", X"EBBB", X"E809", X"2EF0",
		X"92FC", X"92FC", X"E0A1", X"EFBA", X"E404",
		X"2EF0", X"92FC", X"92FC", X"EFAF", X"EFBF",
		X"E809", X"2EF0", X"92FC", X"92FC", X"E0A1",
		X"E0B0", X"E000", X"2EF0", X"92FC", X"92FC",
		X"EFAF", X"E0BF", X"E211", X"931C", X"931C",
		X"910C", X"910C", X"9300", X"0900", X"0900",
		X"E41A", X"9310", X"0FFF", X"0FFF", X"910C",
		X"910C", X"9300", X"0900", X"0900", X"E010",
		X"931C", X"931C", X"910C", X"910C", X"9300",
		X"0900", X"0900", X"EAA0", X"E1B1", X"E302",
		X"2EF0", X"92FD", X"92FD", X"ED0A", X"2EF0",
		X"92FD", X"92FD", X"EFAF", X"EFBF", X"E506",
		X"2EF0", X"92FD", X"92FD", X"E007", X"2EF0",
		X"92FD", X"92FD", X"EBA6", X"E0BA", X"E211",
		X"931C", X"931C", X"910D", X"910D", X"9300",
		X"0900", X"0900", X"E41A", X"9310", X"0AB7",
		X"0AB7", X"910D", X"910D", X"9300", X"0900",
		X"0900", X"E010", X"9310", X"0AB8", X"0AB8",
		X"910D", X"910D", X"9300", X"0900", X"0900",
		X"EAA0", X"E1B1", X"E001", X"2EF0", X"92FE",
		X"92FE", X"E403", X"2EF0", X"92FE", X"92FE",
		X"E0A0", X"E0B0", X"E10F", X"2EF0", X"92FE",
		X"92FE", X"E706", X"2EF0", X"92FE", X"92FE",
		X"E0A9", X"E0BF", X"E211", X"931D", X"931D",
		X"910E", X"910E", X"9300", X"0900", X"0900",
		X"E21B", X"9310", X"0F08", X"0F08", X"910E",
		X"910E", X"9300", X"0900", X"0900", X"E013",
		X"9310", X"0F07", X"0F07", X"910E", X"910E",
		X"9300", X"0900", X"0900", X"EAC0", X"E1D1",
		X"E302", X"2EF0", X"92F9", X"92F9", X"ED0A",
		X"2EF0", X"92F9", X"92F9", X"EFCF", X"EFDF",
		X"E506", X"2EF0", X"92F9", X"92F9", X"E007",
		X"2EF0", X"92F9", X"92F9", X"EAC0", X"E1D1",
		X"E001", X"2EF0", X"92FA", X"92FA", X"E403",
		X"2EF0", X"92FA", X"92FA", X"E0C0", X"E0D0",
		X"E10F", X"2EF0", X"92FA", X"92FA", X"E706",
		X"2EF0", X"92FA", X"92FA", X"E3C3", X"E0D0",
		X"E40D", X"2EF0", X"82FC", X"82FC", X"EE0A",
		X"2EF0", X"8AFF", X"8AFF", X"EACE", X"EFD0",
		X"E30E", X"2EF0", X"AEF9", X"AEF9", X"E60B",
		X"2EF0", X"AEFF", X"AEFF", X"EAE0", X"E1F1",
		X"E302", X"2EF0", X"92F1", X"92F1", X"ED0A",
		X"2EF0", X"92F1", X"92F1", X"EFEF", X"EFFF",
		X"E506", X"2EF0", X"92F1", X"92F1", X"E007",
		X"2EF0", X"92F1", X"92F1", X"EAE0", X"E1F1",
		X"E001", X"2EF0", X"92F2", X"92F2", X"E403",
		X"2EF0", X"92F2", X"92F2", X"E0E0", X"E0F0",
		X"E10F", X"2EF0", X"92F2", X"92F2", X"E706",
		X"2EF0", X"92F2", X"92F2", X"E3E3", X"E0F0",
		X"E40D", X"2EF0", X"82F4", X"82F4", X"EE0A",
		X"2EF0", X"8AF7", X"8AF7", X"EAEE", X"EFF0",
		X"E30E", X"2EF0", X"AEF1", X"AEF1", X"E60B",
		X"2EF0", X"AEF7", X"AEF7", X"E617", X"931F",
		X"931F", X"910F", X"910F", X"9300", X"1000",
		X"1000", X"E810", X"EA25", X"E83F", X"931F",
		X"931F", X"932F", X"932F", X"933F", X"933F",
		X"910F", X"910F", X"90FF", X"90FF", X"90EF",
		X"90EF", X"9300", X"1000", X"1000", X"92F0",
		X"1000", X"1000", X"92E0", X"1000", X"1000",
		X"EA15", X"FD12", X"0000", X"9310", X"1000", X"1000", -- SBRC bubble inserted
		X"FD16", X"0000", X"9310", X"0900", X"E014", X"FD12", X"0000", -- SBRC bubble inserted (x2)
		X"9310", X"1000", X"1000", X"FD14", X"0000", X"9310", -- SBRC bubble inserted
		X"0900", X"E915", X"FD17", X"0000", X"9310", X"1000", -- SBRC bubble inserted
		X"1000", X"FD15", X"0000", X"9310", X"0900", X"E616", -- SBRC bubble inserted
		X"FF15", X"0000", X"9310", X"1000", X"FF10", X"0000", X"9310", -- SBRS bubble inserted (x2)
		X"0900", X"0900", X"EB1E", X"FF14", X"0000", X"9310", -- SBRS bubble inserted
		X"1000", X"FF16", X"0000", X"9310", X"0900", X"0900", -- SBRS bubble inserted
		X"E011", X"FF10", X"0000", X"9310", X"1000", X"FF16", X"0000", -- SBRS bubble inserted (x2)
		X"9310", X"0900", X"0900", X"E000", X"E010",
		X"1301", X"0000", X"9300", X"1000", X"EF0F", X"1301", X"0000", -- CPSE bubble inserted (x2)
		X"9300", X"1000", X"1000", X"EF1F", X"1301", X"0000", -- CPSE bubble inserted 
		X"9310", X"1000", X"1301", X"0000", X"E010", X"E307", -- CPSE bubble inserted 
		X"1301", X"0000", X"9300", X"1000", X"1000", X"E505", -- CPSE bubble inserted
		X"940C", X"1100", X"1100", X"9300", X"1000",
		X"1000", X"E20C", X"940C", X"1134", X"1134",
		X"9300", X"1000", X"1000", X"E404", X"C0C8",
		X"C0C8", X"9300", X"1000", X"1000", X"E001",
		X"C0FC", X"C0FC", X"9300", X"1000", X"1000",
		X"E9E5", X"E1F4", X"E909", X"9409", X"9409",
		X"9300", X"1000", X"1000", X"EDEC", X"E1F4",
		X"E200", X"9409", X"9409", X"9300", X"1000",
		X"1000", X"E80E", X"940E", X"155F", X"155F",
		X"155F", X"9300", X"1000", X"1000", X"9508",
		X"9508", X"9508", X"9508", X"9300", X"0900",
		X"0900", X"E202", X"940E", X"1582", X"1582",
		X"1582", X"9300", X"1000", X"1000", X"9508",
		X"9508", X"9508", X"9508", X"9300", X"0900",
		X"0900", X"E405", X"D178", X"D178", X"D178",
		X"9300", X"1000", X"1000", X"9508", X"9508",
		X"9508", X"9508", X"9300", X"0900", X"0900",
		X"EE0A", X"D216", X"D216", X"D216", X"9300",
		X"1000", X"1000", X"9508", X"9508", X"9508",
		X"9508", X"9300", X"0900", X"0900", X"E007",
		X"EFEF", X"E1F7", X"9509", X"9509", X"9509",
		X"9300", X"1000", X"1000", X"9508", X"9508",
		X"9508", X"9508", X"9300", X"0900", X"0900",
		X"E101", X"E2E2", X"E1F9", X"9509", X"9509",
		X"9509", X"9300", X"1000", X"1000", X"9508",
		X"9508", X"9508", X"9508", X"9300", X"0900",
		X"0900", X"C523", X"C523", X"E909", X"94F8", X"0000", X"0000", X"0000", -- BCLR bubble inserted (x3)
		X"940E", X"1A30", X"1A30", X"1A30", X"9518",
		X"9518", X"9518", X"9518", X"F06F", X"F06F",
		X"E010", X"9300", X"0900", X"0900", X"EE00",
		X"94F8", X"0000", X"0000", X"0000", X"940E", X"1A50", X"1A50", X"1A50", -- BCLR bubble inserted (x3)
		X"9518", X"9518", X"9518", X"9518", X"F0C7",
		X"F0C7", X"E011", X"9300", X"0900", X"0900",
		X"940C", X"1B00", X"1B00", X"EF0F", X"2E00",
		X"920F", X"920F", X"0000", X"901F", X"901F",
		X"1001", X"0000", X"9200", X"1000", X"E001", X"2E10", -- CPSE bubble inserted
		X"921F", X"921F", X"0000", X"902F", X"902F",
		X"1012", X"0000", X"9210", X"1000", X"E002", X"2E20", -- CPSE bubble inserted
		X"922F", X"922F", X"0000", X"903F", X"903F",
		X"1023", X"0000", X"9220", X"1000", X"E003", X"2E30", -- CPSE bubble inserted
		X"923F", X"923F", X"0000", X"904F", X"904F",
		X"1034", X"0000", X"9230", X"1000", X"E004", X"2E40", -- CPSE bubble inserted
		X"924F", X"924F", X"0000", X"905F", X"905F",
		X"1045", X"0000", X"9240", X"1000", X"E005", X"2E50", -- CPSE bubble inserted
		X"925F", X"925F", X"0000", X"906F", X"906F",
		X"1056", X"0000", X"9250", X"1000", X"E006", X"2E60", -- CPSE bubble inserted
		X"926F", X"926F", X"0000", X"907F", X"907F",
		X"1067", X"0000", X"9260", X"1000", X"E007", X"2E70", -- CPSE bubble inserted
		X"927F", X"927F", X"0000", X"908F", X"908F",
		X"1078", X"0000", X"9270", X"1000", X"E008", X"2E80", -- CPSE bubble inserted
		X"928F", X"928F", X"0000", X"909F", X"909F",
		X"1089", X"0000", X"9280", X"1000", X"E009", X"2E90", -- CPSE bubble inserted
		X"929F", X"929F", X"0000", X"90AF", X"90AF",
		X"109A", X"0000", X"9290", X"1000", X"E100", X"2EA0", -- CPSE bubble inserted
		X"92AF", X"92AF", X"0000", X"90BF", X"90BF",
		X"10AB", X"0000", X"92A0", X"1000", X"E101", X"2EB0", -- CPSE bubble inserted
		X"92BF", X"92BF", X"0000", X"90CF", X"90CF",
		X"10BC", X"0000", X"92B0", X"1000", X"E102", X"2EC0", -- CPSE bubble inserted
		X"92CF", X"92CF", X"0000", X"90DF", X"90DF",
		X"10CD", X"0000", X"92C0", X"1000", X"E103", X"2ED0", -- CPSE bubble inserted
		X"92DF", X"92DF", X"0000", X"90EF", X"90EF",
		X"10DE", X"0000", X"92D0", X"1000", X"E104", X"2EE0", -- CPSE bubble inserted
		X"92EF", X"92EF", X"0000", X"90FF", X"90FF",
		X"10EF", X"0000", X"92E0", X"1000", X"E105", X"2EF0", -- CPSE bubble inserted
		X"92FF", X"92FF", X"0000", X"910F", X"910F",
		X"12F0", X"0000", X"92F0", X"1000", X"E106", X"930F", -- CPSE bubble inserted
		X"930F", X"0000", X"911F", X"911F", X"1301", X"0000", -- CPSE bubble inserted
		X"9260", X"1000", X"E117", X"931F", X"931F",
		X"0000", X"912F", X"912F", X"1312", X"0000", X"9270", -- CPSE bubble inserted
		X"1000", X"E128", X"932F", X"932F", X"0000",
		X"913F", X"913F", X"1323", X"0000", X"9320", X"1000", -- CPSE bubble inserted
		X"E139", X"933F", X"933F", X"0000", X"914F",
		X"914F", X"1334", X"0000", X"9330", X"1000", X"E240", -- CPSE bubble inserted
		X"934F", X"934F", X"0000", X"915F", X"915F",
		X"1345", X"0000", X"9340", X"1000", X"E251", X"935F", -- CPSE bubble inserted
		X"935F", X"0000", X"916F", X"916F", X"1356", X"0000", -- CPSE bubble inserted
		X"9350", X"1000", X"E262", X"936F", X"936F",
		X"0000", X"917F", X"917F", X"1367", X"0000", X"9360", -- CPSE bubble inserted
		X"1000", X"E273", X"937F", X"937F", X"0000",
		X"918F", X"918F", X"1378", X"0000", X"9370", X"1000", -- CPSE bubble inserted
		X"E284", X"938F", X"938F", X"0000", X"919F",
		X"919F", X"1389", X"0000", X"9380", X"1000", X"E295", -- CPSE bubble inserted
		X"939F", X"939F", X"0000", X"91AF", X"91AF",
		X"139A", X"0000", X"9390", X"1000", X"E2A6", X"93AF", -- CPSE bubble inserted
		X"93AF", X"0000", X"91BF", X"91BF", X"13AB", X"0000", -- CPSE bubble inserted
		X"93A0", X"1000", X"E2B7", X"93BF", X"93BF",
		X"0000", X"91CF", X"91CF", X"13BC", X"0000", X"93B0", -- CPSE bubble inserted
		X"1000", X"E2C8", X"93CF", X"93CF", X"0000",
		X"91DF", X"91DF", X"13CD", X"0000", X"93C0", X"1000", -- CPSE bubble inserted
		X"E2D9", X"93DF", X"93DF", X"0000", X"91EF",
		X"91EF", X"13DE", X"0000", X"93D0", X"1000", X"E3E0", -- CPSE bubble inserted
		X"93EF", X"93EF", X"0000", X"91FF", X"91FF",
		X"13EF", X"0000", X"93E0", X"1000", X"E3F1", X"93FF", -- CPSE bubble inserted
		X"93FF", X"0000", X"901F", X"901F", X"11F1", X"0000", -- CPSE bubble inserted
		X"93F0", X"1000", X"C10F", X"C10F", X"E400",
		X"E51A", X"1F01", X"0000", X"0000", X"0000", X"F415", X"F415", X"F41C", -- ADC bubble inserted (x3)
		X"F41C", X"F01B", X"F01B", X"F022", X"F022",
		X"F409", X"F409", X"F418", X"F418", X"9300",
		X"1000", X"1000", X"E92A", X"1302", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"ED02", X"1F01", X"0000", X"0000", X"0000", X"F475", X"F475", -- ADC bubble inserted (x3)
		X"F41C", X"F41C", X"F41B", X"F41B", X"F41A",
		X"F41A", X"F421", X"F421", X"F018", X"F018",
		X"9300", X"1000", X"1000", X"E22C", X"1302", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"E708", X"1F01", X"0000", X"0000", X"0000", X"F095", -- ADC bubble inserted (x3)
		X"F095", X"F41C", X"F41C", X"F01B", X"F01B",
		X"F01A", X"F01A", X"F421", X"F421", X"F418",
		X"F418", X"9300", X"1000", X"1000", X"ED23",
		X"1302", X"0000", X"9300", X"0900", X"E400", X"E51A", -- CPSE bubble inserted
		X"0F01", X"0000", X"0000", X"0000", X"F42D", X"F42D", X"F41C", X"F41C", -- ADD bubble inserted (x3)
		X"F013", X"F013", X"F09A", X"F09A", X"F421",
		X"F421", X"F418", X"F418", X"9300", X"1000",
		X"1000", X"E92A", X"1302", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"ED02", X"0F01", X"0000", X"0000", X"0000", X"F40D", X"F40D", X"F41C", -- ADD bubble inserted (x3)
		X"F41C", X"F41B", X"F41B", X"F422", X"F422",
		X"F421", X"F421", X"F018", X"F018", X"9300",
		X"1000", X"1000", X"E22C", X"1302", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"E708", X"0F01", X"0000", X"0000", X"0000", X"F00D", X"F00D", -- ADD bubble inserted (x3)
		X"F41C", X"F41C", X"F01B", X"F01B", X"F01A",
		X"F01A", X"F419", X"F419", X"F418", X"F418",
		X"9300", X"1000", X"1000", X"ED22", X"1302", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"E480", X"E59A", X"96CF", 
		X"96CF", X"0000", X"0000", X"0000", X"F424", X"F424", X"F41B", X"F41B", -- ADIW bubble inserted (x3)
		X"F412", X"F412", X"F419", X"F419", X"F420",
		X"F420", X"9380", X"1000", X"1000", X"9390",
		X"0900", X"0900", X"E7AF", X"E5BA", X"138A", X"0000", -- CPSE bubble inserted
		X"9380", X"0900", X"139B", X"0000", X"9390", X"0900", -- CPSE bubble inserted
		X"EFAF", X"EFBF", X"9612", X"9612", X"0000", X"0000", X"0000", X"F414", -- ADIW bubble inserted (x3)
		X"F414", X"F41B", X"F41B", X"F41A", X"F41A",
		X"F421", X"F421", X"F018", X"F018", X"93A0",
		X"1000", X"1000", X"93B0", X"0900", X"0900",
		X"E0C1", X"E0D0", X"13AC", X"0000", X"93A0", X"0900", -- CPSE bubble inserted
		X"13BD", X"0000", X"93B0", X"0900", X"EFCE", X"EFDF", -- CPSE bubble inserted
		X"96EF", X"96EF", X"0000", X"0000", X"0000", X"F44C", X"F44C", X"F41B", -- ADIW bubble inserted (x3)
		X"F41B", X"F41A", X"F41A", X"F411", X"F411",
		X"F018", X"F018", X"93C0", X"1000", X"1000",
		X"93D0", X"0900", X"0900", X"E3ED", X"E0F0",
		X"13CE", X"0000", X"93C0", X"0900", X"13DF", X"0000", X"93D0", -- CPSE bubble inserted (x2)
		X"0900", X"E400", X"E51A", X"2301", X"0000", X"0000", X"0000", X"F41C", -- AND bubble inserted (x3)
		X"F41C", X"F41B", X"F41B", X"F41A", X"F41A",
		X"F421", X"F421", X"9300", X"1000", X"1000",
		X"E420", X"1302", X"0000", X"9300", X"0900", X"ED02", -- CPSE bubble inserted
		X"2301", X"0000", X"0000", X"0000", X"F414", X"F414", X"F423", X"F423", -- AND bubble inserted (x3)
		X"F422", X"F422", X"F419", X"F419", X"9300",
		X"1000", X"1000", X"E522", X"1302", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"E000", X"2301", X"0000", X"0000", X"0000", X"F41C", X"F41C", -- AND bubble inserted (x3)
		X"F41B", X"F41B", X"F412", X"F412", X"F019",
		X"F019", X"9300", X"1000", X"1000", X"E020",
		X"1302", X"0000", X"9300", X"0900", X"E40F", X"7D0D", X"0000", X"0000", X"0000", -- CPSE bubble inserted & ANDI bubble inserted (x3)
		X"F42C", X"F42C", X"F423", X"F423", X"F41A",
		X"F41A", X"F421", X"F421", X"9300", X"1000",
		X"1000", X"E42D", X"1302", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"7B00", X"0000", X"0000", X"0000", X"F42C", X"F42C", X"F413", X"F413", -- ANDI bubble inserted (x3)
		X"F41A", X"F41A", X"F021", X"F021", X"9300",
		X"1000", X"1000", X"E020", X"1302", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"7702", X"0000", X"0000", X"0000", X"F41C", X"F41C", X"F413", -- ANDI bubble inserted (x3)
		X"F413", X"F41A", X"F41A", X"F021", X"F021",
		X"9300", X"1000", X"1000", X"E020", X"1302", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"EB06", X"9505", X"0000", X"0000", X"0000", X"F414", -- ASR bubble inserted (x3)
		X"F414", X"F023", X"F023", X"F01A", X"F01A",
		X"F419", X"F419", X"F410", X"F410", X"9300",
		X"1000", X"1000", X"ED2B", X"1302", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"E509", X"9505", X"0000", X"0000", X"0000", X"F02C", X"F02C", -- ASR bubble inserted (x3)
		X"F01B", X"F01B", X"F412", X"F412", X"F411",
		X"F411", X"F018", X"F018", X"9300", X"1000",
		X"1000", X"E22C", X"1302", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"EF0F", X"9505", X"0000", X"0000", X"0000", X"F014", X"F014", X"F423", -- ASR bubble inserted (x3)
		X"F423", X"F01A", X"F01A", X"F421", X"F421",
		X"F018", X"F018", X"9300", X"1000", X"1000",
		X"EF2F", X"1302", X"0000", X"9300", X"0900", X"9408", -- CPSE bubble inserted
		X"0000", X"0000", X"0000", X"F018", X"F018", X"9488", X"0000", X"0000", X"0000", X"F410", X"F410", -- BSET bubble inserted (x3) & BCLR bubble inserted (x3)
		X"9418", X"0000", X"0000", X"0000", X"F011", X"F011", X"9498", X"0000", X"0000", X"0000", X"F411", -- BSET bubble inserted (x3) & BCLR bubble inserted (x3)
		X"F411", X"9428", X"0000", X"0000", X"0000", X"F01A", X"F01A", X"94A8", X"0000", X"0000", X"0000", -- BSET bubble inserted (x3) & BCLR bubble inserted (x3)
		X"F412", X"F412", X"9438", X"0000", X"0000", X"0000", X"F01B", X"F01B", -- BSET bubble inserted (x3)
		X"94B8", X"0000", X"0000", X"0000", X"F413", X"F413", X"9448", X"0000", X"0000", X"0000", X"F014", -- BCLR bubble inserted (x3) and BSET bubble inserted (X3)
		X"F014", X"94C8", X"0000", X"0000", X"0000", X"F424", X"F424", X"9458", X"0000", X"0000", X"0000", -- BCLR bubble inserted (x3) and BSET bubble inserted (x3)
		X"F015", X"F015", X"94D8", X"0000", X"0000", X"0000", X"F41D", X"F41D", -- BCLR bubble inserted (x3)
		X"9468", X"0000", X"0000", X"0000", X"F016", X"F016", X"94E8", X"0000", X"0000", X"0000", X"F416", -- BSET bubble inserted (x3) and BCLR bubble inserted (x3)
		X"F416", X"9478", X"0000", X"0000", X"0000", X"F017", X"F017", X"94F8", X"0000", X"0000", X"0000", -- BSET bubble inserted (x3) and BCLR bubble inserted (x3)
		X"F41F", X"F41F", X"0000", X"E503", X"FB04", X"0000", X"0000", X"0000", -- BST bubble inserted (x3)
		X"F01E", X"F01E", X"F907", X"0000", X"0000", X"0000", X"ED13", X"1301", -- BLD bubble inserted (x3)
		X"0000", X"9300", X"1000", X"FB05", X"0000", X"0000", X"0000", X"F41E", X"F41E", -- CPSE bubble inserted & BST bubble inserted (x3)
		X"F901", X"0000", X"0000", X"0000", X"ED11", X"1301", X"0000", X"9300", X"1000", -- BLD bubble inserted (x3) & CPSE bubble inserted
		X"E703", X"9500", X"0000", X"0000", X"0000", X"F01C", X"F01C", X"F41B", -- COM bubble inserted (x3)
		X"F41B", X"F01A", X"F01A", X"F419", X"F419",
		X"F018", X"F018", X"9300", X"1000", X"1000",
		X"E81C", X"1301", X"0000", X"9300", X"0900", X"E000", -- CPSE bubble inserted
		X"9500", X"0000", X"0000", X"0000", X"F00C", X"F00C", X"F41B", X"F41B", -- COM bubble inserted (x3)
		X"F01A", X"F01A", X"F419", X"F419", X"F018",
		X"F018", X"9300", X"1000", X"1000", X"EF1F",
		X"1301", X"0000", X"9300", X"0900", X"E505", X"9500", -- CPSE bubble inserted
		X"0000", X"0000", X"0000", X"F014", X"F014", X"F423", X"F423", X"F01A", -- COM bubble inserted (x3)
		X"F01A", X"F419", X"F419", X"F018", X"F018",
		X"9300", X"1000", X"1000", X"EA1A", X"1301", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"E703", X"EF10", X"1701", X"0000", X"0000", X"0000", -- CP bubble inserted (x3)
		X"F41D", X"F41D", X"F41C", X"F41C", X"F023",
		X"F023", X"F01A", X"F01A", X"F411", X"F411",
		X"F010", X"F010", X"9300", X"1000", X"1000",
		X"E004", X"E013", X"1701", X"0000", X"0000", X"0000", X"F425", X"F425", -- CP bubble inserted (x3)
		X"F414", X"F414", X"F413", X"F413", X"F41A",
		X"F41A", X"F419", X"F419", X"F418", X"F418",
		X"9300", X"1000", X"1000", X"E505", X"EA1A",
		X"1701", X"0000", X"0000", X"0000", X"F025", X"F025", X"F41C", X"F41C", -- CP bubble inserted (x3)
		X"F013", X"F013", X"F01A", X"F01A", X"F411",
		X"F411", X"F018", X"F018", X"9300", X"1000",
		X"1000", X"E703", X"EF10", X"9408", X"0000", X"0000", X"0000", X"0701", X"0000", X"0000", X"0000", -- BSET bubble inserted (x3) & CPC bubble inserted (x3)
		X"F41D", X"F41D", X"F41C", X"F41C", X"F01B",
		X"F01B", X"F012", X"F012", X"F411", X"F411",
		X"F018", X"F018", X"9300", X"1000", X"1000",
		X"E004", X"E013", X"9408", X"0000", X"0000", X"0000", X"0701", X"0000", X"0000", X"0000", X"F41D", -- BSET bubble inserted (x3) & CPC bubble inserted (x3)
		X"F41D", X"F414", X"F414", X"F423", X"F423",
		X"F41A", X"F41A", X"F411", X"F411", X"F410",
		X"F410", X"9300", X"1000", X"1000", X"E004",
		X"E013", X"9418", X"0000", X"0000", X"0000", X"9408", X"0000", X"0000", X"0000", X"0701", X"0000", X"0000", X"0000", X"F425", -- x2 BSET bubble inserted (x3) & CPC bubble inserted (x3)
		X"F425", X"F41C", X"F41C", X"F41B", X"F41B",
		X"F41A", X"F41A", X"F019", X"F019", X"F418",
		X"F418", X"9300", X"1000", X"1000", X"E400",
		X"330F", X"0000", X"0000", X"0000", X"F01D", X"F01D", X"F41C", X"F41C", -- CPI bubble inserted (x3)
		X"F41B", X"F41B", X"F41A", X"F41A", X"F419",
		X"F419", X"F418", X"F418", X"9300", X"1000",
		X"1000", X"E008", X"3000", X"0000", X"0000", X"0000", X"F41D", X"F41D", -- CPI bubble inserted (x3)
		X"F41C", X"F41C", X"F41B", X"F41B", X"F41A",
		X"F41A", X"F419", X"F419", X"F418", X"F418",
		X"9300", X"1000", X"1000", X"E901", X"300E", X"0000", X"0000", X"0000", -- CPI bubble inserted (x3)
		X"F02D", X"F02D", X"F01C", X"F01C", X"F41B",
		X"F41B", X"F012", X"F012", X"F419", X"F419",
		X"F418", X"F418", X"9300", X"1000", X"1000",
		X"EF0F", X"950A", X"0000", X"0000", X"0000", X"F01C", X"F01C", X"F41B", -- DEC bubble inserted (x3)
		X"F41B", X"F022", X"F022", X"F419", X"F419",
		X"9300", X"1000", X"1000", X"EF1E", X"1301", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"9503", X"0000", X"0000", X"0000", X"9503", X"0000", X"0000", X"0000", X"F41C", -- x2 INC bubble inserted (x3)
		X"F41C", X"F41B", X"F41B", X"F41A", X"F41A",
		X"F011", X"F011", X"9300", X"1000", X"1000",
		X"E010", X"1301", X"0000", X"9300", X"0900", X"EF06", -- CPSE bubble inserted
		X"E619", X"2701", X"0000", X"0000", X"0000", X"F014", X"F014", X"F41B", -- EOR bubble inserted (x3)
		X"F41B", X"F022", X"F022", X"F419", X"F419",
		X"9300", X"1000", X"1000", X"E91F", X"1301", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"E505", X"EE14", X"2701", X"0000", X"0000", X"0000", -- EOR bubble inserted (x3)
		X"F014", X"F014", X"F41B", X"F41B", X"F012",
		X"F012", X"F419", X"F419", X"9300", X"1000",
		X"1000", X"EB11", X"1301", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"E708", X"EF1F", X"2701", X"0000", X"0000", X"0000", X"F01C", X"F01C", -- EOR bubble inserted (x3)
		X"F413", X"F413", X"F022", X"F022", X"F419",
		X"F419", X"9300", X"1000", X"1000", X"E817",
		X"1301", X"0000", X"9300", X"0900", X"EF06", X"9506", -- CPSE bubble inserted
		X"0000", X"0000", X"0000", X"F41C", X"F41C", X"F41B", X"F41B", X"F412", -- LSR bubble inserted (x3)
		X"F412", X"F419", X"F419", X"F420", X"F420",
		X"9300", X"1000", X"1000", X"E71B", X"1301", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"E505", X"9506", X"0000", X"0000", X"0000", X"F014", -- LSR bubble inserted (x3)
		X"F014", X"F023", X"F023", X"F41A", X"F41A",
		X"F411", X"F411", X"F018", X"F018", X"9300",
		X"1000", X"1000", X"E21A", X"1301", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"E708", X"9506", X"0000", X"0000", X"0000", X"F414", X"F414", -- LSR bubble inserted (x3)
		X"F41B", X"F41B", X"F42A", X"F42A", X"F419",
		X"F419", X"F410", X"F410", X"9300", X"1000",
		X"1000", X"E31C", X"1301", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"EF06", X"9501", X"0000", X"0000", X"0000", X"F424", X"F424", X"F413", -- NEG bubble inserted (x3)
		X"F413", X"F41A", X"F41A", X"F421", X"F421",
		X"F018", X"F018", X"9300", X"1000", X"1000",
		X"E01A", X"1301", X"0000", X"9300", X"0900", X"E505", -- CPSE bubble inserted
		X"9501", X"0000", X"0000", X"0000", X"F01C", X"F01C", X"F41B", X"F41B", -- NEG bubble inserted (x3)
		X"F012", X"F012", X"F419", X"F419", X"F020",
		X"F020", X"9300", X"1000", X"1000", X"EA1B",
		X"1301", X"0000", X"9300", X"0900", X"E708", X"9501", -- CPSE bubble inserted
		X"0000", X"0000", X"0000", X"F02C", X"F02C", X"F41B", X"F41B", X"F01A", -- NEG bubble inserted (x3)
		X"F01A", X"F419", X"F419", X"F028", X"F028",
		X"9300", X"1000", X"1000", X"E818", X"1301", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"EF06", X"E914", X"2B01", X"0000", X"0000", X"0000", -- OR bubble inserted (x3)
		X"F034", X"F034", X"F41B", X"F41B", X"F012",
		X"F012", X"F419", X"F419", X"9300", X"1000",
		X"1000", X"EF16", X"1301", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"E505", X"E71E", X"2B01", X"0000", X"0000", X"0000", X"F424", X"F424", -- OR bubble inserted (x3)
		X"F423", X"F423", X"F41A", X"F41A", X"F419",
		X"F419", X"9300", X"1000", X"1000", X"E71F",
		X"1301", X"0000", X"9300", X"0900", X"E708", X"EF1F", -- CPSE bubble inserted
		X"2B01", X"0000", X"0000", X"0000", X"F024", X"F024", X"F413", X"F413", -- OR bubble inserted (x3)
		X"F012", X"F012", X"F419", X"F419", X"9300",
		X"1000", X"1000", X"EF1F", X"1301", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"EF06", X"6D0D", X"0000", X"0000", X"0000", X"F01C", X"F01C", -- ORI bubble inserted (x3)
		X"F41B", X"F41B", X"F01A", X"F01A", X"F419",
		X"F419", X"9300", X"1000", X"1000", X"EF1F",
		X"1301", X"0000", X"9300", X"0900", X"E505", X"6102", -- CPSE bubble inserted
		X"0000", X"0000", X"0000", X"F41C", X"F41C", X"F41B", X"F41B", X"F41A", -- ORI bubble inserted (x3)
		X"F41A", X"F419", X"F419", X"9300", X"1000",
		X"1000", X"E517", X"1301", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"E708", X"6000", X"0000", X"0000", X"0000", X"F424", X"F424", X"F423", -- ORI bubble inserted (x3)
		X"F423", X"F41A", X"F41A", X"F411", X"F411",
		X"9300", X"1000", X"1000", X"E718", X"1301", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"9488", X"0000", X"0000", X"0000", X"EF06", X"9507", X"0000", X"0000", X"0000", -- BCLR bubble inserted (x3) & ROR bubble inserted (x3)
		X"F41C", X"F41C", X"F413", X"F413", X"F412",
		X"F412", X"F429", X"F429", X"F418", X"F418",
		X"9300", X"1000", X"1000", X"E71B", X"1301", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"E505", X"9507", X"0000", X"0000", X"0000", X"F01C", -- ROR bubble inserted (x3)
		X"F01C", X"F01B", X"F01B", X"F412", X"F412",
		X"F411", X"F411", X"F018", X"F018", X"9300",
		X"1000", X"1000", X"E21A", X"1301", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"E708", X"9507", X"0000", X"0000", X"0000", X"F41C", X"F41C", -- ROR bubble inserted (x3)
		X"F01B", X"F01B", X"F01A", X"F01A", X"F419",
		X"F419", X"F418", X"F418", X"9300", X"1000",
		X"1000", X"EB1C", X"1301", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"9488", X"0000", X"0000", X"0000", X"E400", X"E51A", X"0B01", X"0000", X"0000", X"0000", X"F02D", -- BCLR bubble inserted (x3) & SBC bubble inserted (x3)
		X"F02D", X"F01C", X"F01C", X"F41B", X"F41B",
		X"F01A", X"F01A", X"F419", X"F419", X"F018",
		X"F018", X"9300", X"1000", X"1000", X"EE26",
		X"1302", X"0000", X"9300", X"0900", X"ED02", X"0B01", X"0000", X"0000", X"0000", -- CPSE bubble inserted & SBC bubble inserted (x3)
		X"F01D", X"F01D", X"F01C", X"F01C", X"F01B",
		X"F01B", X"F41A", X"F41A", X"F419", X"F419",
		X"F418", X"F418", X"9300", X"1000", X"1000",
		X"E727", X"1302", X"0000", X"9300", X"0900", X"E708", -- CPSE bubble inserted
		X"0B01", X"0000", X"0000", X"0000", X"F01D", X"F01D", X"F41C", X"F41C", -- SBC bubble inserted (x3)
		X"F41B", X"F41B", X"F41A", X"F41A", X"F419",
		X"F419", X"F418", X"F418", X"9300", X"1000",
		X"1000", X"E12E", X"1302", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"9488", X"0000", X"0000", X"0000", X"E400", X"4606", X"0000", X"0000", X"0000", X"F035", X"F035", -- BCLR bubble inserted (x3) and SBCI bubble inserted (x3)
		X"F01C", X"F01C", X"F41B", X"F41B", X"F01A",
		X"F01A", X"F419", X"F419", X"F018", X"F018",
		X"9300", X"1000", X"1000", X"ED2A", X"1302", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"ED02", X"4203", X"0000", X"0000", X"0000", X"F02D", -- SBCI bubble inserted (x3)
		X"F02D", X"F01C", X"F01C", X"F413", X"F413",
		X"F012", X"F012", X"F419", X"F419", X"F418",
		X"F418", X"9300", X"1000", X"1000", X"EA2E",
		X"1302", X"0000", X"9300", X"0900", X"E708", X"4F0F", X"0000", X"0000", X"0000", -- CPSE bubble inserted & SBCI bubble inserted (x3)
		X"F02D", X"F02D", X"F41C", X"F41C", X"F413",
		X"F413", X"F412", X"F412", X"F419", X"F419",
		X"F018", X"F018", X"9300", X"1000", X"1000",
		X"E729", X"1302", X"0000", X"9300", X"0900", X"E480", -- CPSE bubble inserted
		X"E59A", X"97CF", X"97CF", X"0000", X"0000", X"0000", X"F424", X"F424", -- SBIW bubble inserted (x3)
		X"F41B", X"F41B", X"F412", X"F412", X"F411",
		X"F411", X"F418", X"F418", X"9380", X"1000",
		X"1000", X"9390", X"0900", X"0900", X"E0A1",
		X"E5BA", X"138A", X"0000", X"9380", X"0900", X"139B", X"0000", -- x2 CPSE bubble inserted
		X"9390", X"0900", X"EFAF", X"EFBF", X"9712",
		X"9712", X"0000", X"0000", X"0000", X"F024", X"F024", X"F41B", X"F41B", -- SBIW bubble inserted (x3)
		X"F01A", X"F01A", X"F419", X"F419", X"F418",
		X"F418", X"93A0", X"1000", X"1000", X"93B0",
		X"0900", X"0900", X"EFCD", X"EFDF", X"13AC", X"0000", -- CPSE bubble inserted
		X"93A0", X"0900", X"13BD", X"0000", X"93B0", X"0900", -- CPSE bubble inserted
		X"E0C0", X"E0D0", X"97EF", X"97EF", X"0000", X"0000", X"0000", X"F024", -- SBIW bubble inserted
		X"F024", X"F41B", X"F41B", X"F01A", X"F01A",
		X"F419", X"F419", X"F018", X"F018", X"93C0",
		X"1000", X"1000", X"93D0", X"0900", X"0900",
		X"ECE1", X"EFFF", X"13CE", X"0000", X"93C0", X"0900", -- CPSE bubble inserted
		X"13DF", X"0000", X"93D0", X"0900", X"E400", X"E51A", -- CPSE bubble inserted
		X"1B01", X"0000", X"0000", X"0000", X"F025", X"F025", X"F01C", X"F01C", -- SUB bubble inserted (x3)
		X"F41B", X"F41B", X"F01A", X"F01A", X"F419",
		X"F419", X"F018", X"F018", X"9300", X"1000",
		X"1000", X"EE26", X"1302", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"ED02", X"1B01", X"0000", X"0000", X"0000", X"F01D", X"F01D", X"F01C", -- SUB bubble inserted (x3)
		X"F01C", X"F01B", X"F01B", X"F49A", X"F49A",
		X"F419", X"F419", X"F418", X"F418", X"9300",
		X"1000", X"1000", X"E728", X"1302", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"E708", X"1B01", X"0000", X"0000", X"0000", X"F01D", X"F01D", -- SUB bubble inserted (x3)
		X"F41C", X"F41C", X"F41B", X"F41B", X"F41A",
		X"F41A", X"F419", X"F419", X"F418", X"F418",
		X"9300", X"1000", X"1000", X"E12E", X"1302", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"E400", X"5F0F", X"0000", X"0000", X"0000", X"F01D", -- SUBI bubble inserted (x3)
		X"F01D", X"F41C", X"F41C", X"F41B", X"F41B",
		X"F41A", X"F41A", X"F419", X"F419", X"F018",
		X"F018", X"9300", X"1000", X"1000", X"E421",
		X"1302", X"0000", X"9300", X"0900", X"ED02", X"5707", -- CPSE bubble inserted
		X"0000", X"0000", X"0000", X"F01D", X"F01D", X"F01C", X"F01C", X"F01B", -- SUBI bubble inserted (x3)
		X"F01B", X"F41A", X"F41A", X"F419", X"F419",
		X"F418", X"F418", X"9300", X"1000", X"1000",
		X"E52B", X"1302", X"0000", X"9300", X"0900", X"E708", -- CPSE bubble inserted
		X"5000", X"0000", X"0000", X"0000", X"F41D", X"F41D", X"F41C", X"F41C", -- SUBI bubble inserted (x3)
		X"F41B", X"F41B", X"F41A", X"F41A", X"F419",
		X"F419", X"F418", X"F418", X"9300", X"1000",
		X"1000", X"E728", X"1302", X"0000", X"9300", X"0900", -- CPSE bubble inserted
		X"E10E", X"EE11", X"9502", X"1301", X"0000", X"9300", -- CPSE bubble inserted
		X"0900", X"E00F", X"EF10", X"9502", X"1301", X"0000", -- CPSE bubble inserted
		X"9300", X"0900", X"E101", X"E111", X"9502",
		X"1301", X"0000", X"9300", X"0900", X"E30C", X"E813", -- CPSE bubble inserted
		X"9F01", X"9F01", X"0000", X"0000", X"0000", X"F511", X"F511", X"F418", -- MUL bubble inserted (x3)
		X"F418", X"EB24", X"E13E", X"1120", X"0000", X"9200", -- CPSE bubble inserted
		X"0900", X"1131", X"0000", X"9210", X"0900", X"EF04", -- CPSE bubble inserted
		X"E010", X"9F01", X"9F01", X"0000", X"0000", X"0000", X"F081", X"F081", -- MUL bubble inserted (x3)
		X"F418", X"F418", X"E020", X"E030", X"1120", X"0000", -- CPSE bubble inserted
		X"9200", X"0900", X"1131", X"0000", X"9210", X"0900", -- CPSE bubble inserted
		X"EF0F", X"EF1F", X"9F01", X"9F01", X"0000", X"0000", X"0000", X"F481", -- MUL bubble inserted (x3)
		X"F481", X"F018", X"F018", X"E021", X"EF3E",
		X"1120", X"0000", X"9200", X"0900", X"1131", X"0000", X"9210", -- x2 CPSE bubble inserted 
		X"0900", X"0000", X"0000", X"0000" -- ending buffer
		);

	-- Program Address Bus Test Vector
	constant ProgABTest : testarray := (
		"----------------", "----------------", "----------------", X"0000",            X"0001",            X"0002",            "----------------", X"0003",
		X"0004",            X"0005",            "----------------", X"0006",            X"0007",
		X"0008",            "----------------", X"0009",            X"000A",            X"000B",
		"----------------", X"000C",            X"000D",            X"000E",            "----------------",
		X"000F",            X"0010",            "----------------", X"0011",            X"0012",
		"----------------", X"0013",            X"0014",            X"0015",            "----------------",
		X"0016",            X"0017",            "----------------", X"0018",            X"0019",
		"----------------", X"001A",            X"001B",            X"001C",            "----------------",
		X"001D",            X"001E",            "----------------", X"001F",            X"0020",
		"----------------", X"0021",            X"0022",            X"0023",            "----------------",
		X"0024",            X"0025",            "----------------", X"0026",            X"0027",
		"----------------", X"0028",            X"0029",            X"002A",            X"002B",
		"----------------", X"002C",            X"002D",            X"002E",            X"002F",
		"----------------", X"0030",            X"0031",            X"0032",            X"0033",
		"----------------", X"0034",            X"0035",            X"0036",            X"0037",
		"----------------", X"0038",            X"0039",            X"003A",            X"003B",
		X"003C",            "----------------", X"003D",            X"003E",            X"003F",
		X"0040",            X"0041",            "----------------", X"0042",            X"0043",
		X"0044",            X"0045",            X"0046",            "----------------", X"0047",
		X"0048",            X"0049",            X"004A",            X"004B",            "----------------",
		X"004C",            X"004D",            X"004E",            X"004F",            "----------------",
		X"0050",            "----------------", X"0051",            X"0052",            "----------------",
		X"0053",            X"0054",            X"0055",            "----------------", X"0056",
		"----------------", X"0057",            X"0058",            "----------------", X"0059",
		X"005A",            "----------------", X"005B",            "----------------", X"005C",
		X"005D",            "----------------", X"005E",            X"005F",            X"0060",
		X"0061",            X"0062",            "----------------", X"0063",            X"0064",
		X"0065",            "----------------", X"0066",            X"0067",            X"0068",
		X"0069",            X"006A",            "----------------", X"006B",            X"006C",
		X"006D",            "----------------", X"006E",            X"006F",            X"0070",
		X"0071",            "----------------", X"0072",            "----------------", X"0073",
		X"0074",            "----------------", X"0075",            X"0076",            X"0077",
		"----------------", X"0078",            "----------------", X"0079",            X"007A",
		"----------------", X"007B",            X"007C",            X"007D",            "----------------",
		X"007E",            "----------------", X"007F",            X"0080",            "----------------",
		X"0081",            X"0082",            X"0083",            X"0084",            X"0085",
		"----------------", X"0086",            X"0087",            X"0088",            "----------------",
		X"0089",            X"008A",            X"008B",            X"008C",            X"008D",
		"----------------", X"008E",            X"008F",            X"0090",            "----------------",
		X"0091",            X"0092",            X"0093",            X"0094",            "----------------",
		X"0095",            "----------------", X"0096",            X"0097",            "----------------",
		X"0098",            X"0099",            X"009A",            "----------------", X"009B",
		"----------------", X"009C",            X"009D",            "----------------", X"009E",
		X"009F",            X"00A0",            "----------------", X"00A1",            "----------------",
		X"00A2",            X"00A3",            "----------------", X"00A4",            X"00A5",
		X"00A6",            X"00A7",            X"00A8",            "----------------", X"00A9",
		X"00AA",            X"00AB",            "----------------", X"00AC",            X"00AD",
		X"00AE",            X"00AF",            X"00B0",            "----------------", X"00B1",
		X"00B2",            X"00B3",            "----------------", X"00B4",            X"00B5",
		X"00B6",            X"00B7",            X"00B8",            "----------------", X"00B9",
		X"00BA",            X"00BB",            "----------------", X"00BC",            X"00BD",
		X"00BE",            X"00BF",            X"00C0",            "----------------", X"00C1",
		X"00C2",            X"00C3",            "----------------", X"00C4",            X"00C5",
		X"00C6",            X"00C7",            X"00C8",            "----------------", X"00C9",
		X"00CA",            X"00CB",            "----------------", X"00CC",            X"00CD",
		X"00CE",            X"00CF",            X"00D0",            "----------------", X"00D1",
		X"00D2",            X"00D3",            "----------------", X"00D4",            X"00D5",
		X"00D6",            X"00D7",            X"00D8",            "----------------", X"00D9",
		X"00DA",            X"00DB",            "----------------", X"00DC",            X"00DD",
		X"00DE",            X"00DF",            X"00E0",            "----------------", X"00E1",
		X"00E2",            X"00E3",            "----------------", X"00E4",            X"00E5",
		X"00E6",            X"00E7",            X"00E8",            "----------------", X"00E9",
		X"00EA",            X"00EB",            "----------------", X"00EC",            X"00ED",
		X"00EE",            X"00EF",            X"00F0",            "----------------", X"00F1",
		X"00F2",            X"00F3",            "----------------", X"00F4",            X"00F5",
		X"00F6",            X"00F7",            X"00F8",            "----------------", X"00F9",
		X"00FA",            X"00FB",            "----------------", X"00FC",            X"00FD",
		X"00FE",            X"00FF",            X"0100",            "----------------", X"0101",
		X"0102",            X"0103",            "----------------", X"0104",            X"0105",
		"----------------", X"0106",            "----------------", X"0107",            X"0108",
		"----------------", X"0109",            X"010A",            X"010B",            X"010C",
		"----------------", X"010D",            "----------------", X"010E",            "----------------",
		X"010F",            "----------------", X"0110",            "----------------", X"0111",
		"----------------", X"0112",            X"0113",            "----------------", X"0114",
		X"0115",            "----------------", X"0116",            X"0117",            "----------------",
		X"0118",            X"0119",            "----------------", X"011A",            X"011B",            "----------------", -- SBRC bubble inserted
		X"011C",            "----------------", X"011D",            X"011E",            X"011F",            X"0120", "----------------", -- SBRC bubble inserted (x2)
		X"0121",            X"0122",            "----------------", X"0123",            "----------------", X"0124", -- SBRC bubble inserted
		X"0125",            X"0126",            X"0127",            "----------------", X"0128",            X"0129", -- SBRC bubble inserted
		"----------------", X"012A",            "----------------", X"012B",            X"012C",            X"012D", -- SBRC bubble inserted
		X"012E",            "----------------", X"012F",            X"0130",            X"0131",            "----------------", X"0132", -- SBRS bubble inserted (x2)
		X"0133",            "----------------", X"0134",            X"0135",            "----------------", X"0136", -- SBRS bubble inserted
		X"0137",            X"0138",            "----------------", X"0139",            X"013A",            "----------------", -- SBRS bubble inserted
		X"013B",            X"013C",            "----------------", X"013D",            X"013E",            X"013F", "----------------", -- SBRS bubble inserted (x2)
		X"0140",            X"0141",            "----------------", X"0142",            X"0143",
		X"0144",            "----------------", X"0145",            X"0146",            X"0147",            X"0148", "----------------", -- CPSE bubble inserted (x2)
		X"0149",            X"014A",            "----------------", X"014B",            X"014C", "----------------", -- CPSE bubble inserted
		X"014D",            X"014E",            X"014F",            "----------------", X"0150",            X"0151", -- CPSE bubble inserted
		X"0152",            "----------------", X"0153",            X"0154",            "----------------", X"0155", -- CPSE bubble inserted
		X"0156",            X"0157",            "----------------", X"1100",            X"1101",
		"----------------", X"1102",            X"1103",            X"1104",            "----------------",
		X"1134",            X"1135",            "----------------", X"1136",            X"1137",
		"----------------", X"1200",            X"1201",            "----------------", X"1202",
		X"1203",            "----------------", X"1300",            X"1301",            "----------------",
		X"1302",            X"1303",            X"1304",            X"1305",            "----------------",
		X"1495",            X"1496",            "----------------", X"1497",            X"1498",
		X"1499",            X"149A",            "----------------", X"14DC",            X"14DD",
		"----------------", X"14DE",            X"14DF",            X"14E0",            "----------------",
		"----------------", X"155F",            X"1560",            "----------------", X"1561",
		"----------------", "----------------", "----------------", X"14E1",            X"14E2",
		"----------------", X"14E3",            X"14E4",            X"14E5",            "----------------",
		"----------------", X"1582",            X"1583",            "----------------", X"1584",
		"----------------", "----------------", "----------------", X"14E6",            X"14E7",
		"----------------", X"14E8",            X"14E9",            "----------------", "----------------",
		X"1662",            X"1663",            "----------------", X"1664",            "----------------",
		"----------------", "----------------", X"14EA",            X"14EB",            "----------------",
		X"14EC",            X"14ED",            "----------------", "----------------", X"1704",
		X"1705",            "----------------", X"1706",            "----------------", "----------------",
		"----------------", X"14EE",            X"14EF",            "----------------", X"14F0",
		X"14F1",            X"14F2",            X"14F3",            "----------------", "----------------",
		X"17FF",            X"1800",            "----------------", X"1801",            "----------------",
		"----------------", "----------------", X"14F4",            X"14F5",            "----------------",
		X"14F6",            X"14F7",            X"14F8",            X"14F9",            "----------------",
		"----------------", X"1922",            X"1923",            "----------------", X"1924",
		"----------------", "----------------", "----------------", X"14FA",            X"14FB",
		"----------------", X"14FC",            "----------------", X"1A20",            X"1A21",            "----------------", "----------------", "----------------", -- BCLR bubble inserted (x3)
		X"1A22",            X"1A23",            "----------------", "----------------", X"1A30",
		"----------------", "----------------", "----------------", X"1A24",            "----------------",
		X"1A32",            X"1A33",            X"1A34",            "----------------", X"1A35",
		X"1A36",            "----------------", "----------------", "----------------", X"1A37",            X"1A38",            "----------------", "----------------", -- BCLR bubble inserted (x3)
		X"1A50",            "----------------", "----------------", "----------------", X"1A39",
		"----------------", X"1A52",            X"1A53",            X"1A54",            "----------------",
		X"1A55",            X"1A56",            "----------------", X"1B00",            X"1B01",
		X"1B02",            "----------------", X"1B03",            X"1B04",            "----------------",
		X"1B05",            "----------------", X"1B06",            X"1B07",            X"1B08",            X"1B09", -- CPSE bubble inserted
		X"1B0A",            "----------------", X"1B0B",            X"1B0C",            "----------------",
		X"1B0D",            "----------------", X"1B0E",            X"1B0F",            X"1B10",            X"1B11", -- CPSE bubble inserted
		X"1B12",            "----------------", X"1B13",            X"1B14",            "----------------",
		X"1B15",            "----------------", X"1B16",            X"1B17",            X"1B18",            X"1B19", -- CPSE bubble inserted
		X"1B1A",            "----------------", X"1B1B",            X"1B1C",            "----------------",
		X"1B1D",            "----------------", X"1B1E",            X"1B1F",            X"1B20",            X"1B21", -- CPSE bubble inserted
		X"1B22",            "----------------", X"1B23",            X"1B24",            "----------------",
		X"1B25",            "----------------", X"1B26",            X"1B27",            X"1B28",            X"1B29", -- CPSE bubble inserted
		X"1B2A",            "----------------", X"1B2B",            X"1B2C",            "----------------",
		X"1B2D",            "----------------", X"1B2E",            X"1B2F",            X"1B30",            X"1B31", -- CPSE bubble inserted
		X"1B32",            "----------------", X"1B33",            X"1B34",            "----------------",
		X"1B35",            "----------------", X"1B36",            X"1B37",            X"1B38",            X"1B39", -- CPSE bubble inserted
		X"1B3A",            "----------------", X"1B3B",            X"1B3C",            "----------------",
		X"1B3D",            "----------------", X"1B3E",            X"1B3F",            X"1B40",            X"1B41", -- CPSE bubble inserted
		X"1B42",            "----------------", X"1B43",            X"1B44",            "----------------",
		X"1B45",            "----------------", X"1B46",            X"1B47",            X"1B48",            X"1B49", -- CPSE bubble inserted
		X"1B4A",            "----------------", X"1B4B",            X"1B4C",            "----------------",
		X"1B4D",            "----------------", X"1B4E",            X"1B4F",            X"1B50",            X"1B51", -- CPSE bubble inserted
		X"1B52",            "----------------", X"1B53",            X"1B54",            "----------------",
		X"1B55",            "----------------", X"1B56",            X"1B57",            X"1B58",            X"1B59", -- CPSE bubble inserted
		X"1B5A",            "----------------", X"1B5B",            X"1B5C",            "----------------",
		X"1B5D",            "----------------", X"1B5E",            X"1B5F",            X"1B60",            X"1B61", -- CPSE bubble inserted
		X"1B62",            "----------------", X"1B63",            X"1B64",            "----------------",
		X"1B65",            "----------------", X"1B66",            X"1B67",            X"1B68",            X"1B69", -- CPSE bubble inserted
		X"1B6A",            "----------------", X"1B6B",            X"1B6C",            "----------------",
		X"1B6D",            "----------------", X"1B6E",            X"1B6F",            X"1B70",            X"1B71", -- CPSE bubble inserted
		X"1B72",            "----------------", X"1B73",            X"1B74",            "----------------",
		X"1B75",            "----------------", X"1B76",            X"1B77",            X"1B78",            X"1B79", -- CPSE bubble inserted
		X"1B7A",            "----------------", X"1B7B",            X"1B7C",            "----------------",
		X"1B7D",            "----------------", X"1B7E",            X"1B7F",            X"1B80",            X"1B81", -- CPSE bubble inserted
		"----------------", X"1B82",            X"1B83",            "----------------", X"1B84",            "----------------", -- CPSE bubble inserted
		X"1B85",            X"1B86",            X"1B87",            X"1B88",            "----------------",
		X"1B89",            X"1B8A",            "----------------", X"1B8B",            "----------------", X"1B8C", -- CPSE bubble inserted
		X"1B8D",            X"1B8E",            X"1B8F",            "----------------", X"1B90",
		X"1B91",            "----------------", X"1B92",            "----------------", X"1B93",            X"1B94", -- CPSE bubble inserted
		X"1B95",            X"1B96",            "----------------", X"1B97",            X"1B98",
		"----------------", X"1B99",            "----------------", X"1B9A",            X"1B9B",            X"1B9C", -- CPSE bubble inserted
		X"1B9D",            "----------------", X"1B9E",            X"1B9F",            "----------------",
		X"1BA0",            "----------------", X"1BA1",            X"1BA2",            X"1BA3",            X"1BA4", -- CPSE bubble inserted
		"----------------", X"1BA5",            X"1BA6",            "----------------", X"1BA7",            "----------------", -- CPSE bubble inserted
		X"1BA8",            X"1BA9",            X"1BAA",            X"1BAB",            "----------------",
		X"1BAC",            X"1BAD",            "----------------", X"1BAE",            "----------------", X"1BAF", -- CPSE bubble inserted
		X"1BB0",            X"1BB1",            X"1BB2",            "----------------", X"1BB3",
		X"1BB4",            "----------------", X"1BB5",            "----------------", X"1BB6",            X"1BB7", -- CPSE bubble inserted
		X"1BB8",            X"1BB9",            "----------------", X"1BBA",            X"1BBB",
		"----------------", X"1BBC",            "----------------", X"1BBD",            X"1BBE",            X"1BBF", -- CPSE bubble inserted
		X"1BC0",            "----------------", X"1BC1",            X"1BC2",            "----------------",
		X"1BC3",            "----------------", X"1BC4",            X"1BC5",            X"1BC6",            X"1BC7", -- CPSE bubble inserted
		"----------------", X"1BC8",            X"1BC9",            "----------------", X"1BCA",            "----------------", -- CPSE bubble inserted
		X"1BCB",            X"1BCC",            X"1BCD",            X"1BCE",            "----------------",
		X"1BCF",            X"1BD0",            "----------------", X"1BD1",            "----------------", X"1BD2", -- CPSE bubble inserted
		X"1BD3",            X"1BD4",            X"1BD5",            "----------------", X"1BD6",
		X"1BD7",            "----------------", X"1BD8",            "----------------", X"1BD9",            X"1BDA", -- CPSE bubble inserted
		X"1BDB",            X"1BDC",            "----------------", X"1BDD",            X"1BDE",
		"----------------", X"1BDF",            "----------------", X"1BE0",            X"1BE1",            X"1BE2", -- CPSE bubble inserted
		X"1BE3",            "----------------", X"1BE4",            X"1BE5",            "----------------",
		X"1BE6",            "----------------", X"1BE7",            X"1BE8",            X"1BE9",            X"1BEA", -- CPSE bubble inserted
		"----------------", X"1BEB",            X"1BEC",            "----------------", X"1BED",           "----------------", -- CPSE bubble inserted
		X"1BEE",            X"1BEF",            X"1BF0",            "----------------", X"1D00",
		X"1D01",            X"1D02",            "----------------", "----------------", "----------------", X"1D03",            "----------------", X"1D06", -- ADC bubble inserted (x3)
		"----------------", X"1D0A",            "----------------", X"1D0E",            "----------------",
		X"1D13",            "----------------", X"1D15",            "----------------", X"1D19",
		X"1D1A",            "----------------", X"1D1B",            X"1D1C",            "----------------", X"1D1D", -- CPSE bubble inserted
		X"1D1E",            X"1D1F",            X"1D20",            "----------------", "----------------", "----------------", X"1D21",            "----------------", -- ADC bubble inserted (x3)
		X"1D30",            "----------------", X"1D34",            "----------------", X"1D38",
		"----------------", X"1D3C",            "----------------", X"1D41",            "----------------",
		X"1D45",            X"1D46",            "----------------", X"1D47",            X"1D48",            "----------------",  -- CPSE bubble inserted
		X"1D49",            X"1D4A",            X"1D4B",            X"1D4C",            "----------------", "----------------", "----------------", X"1D4D", -- ADC bubble inserted (x3)
		"----------------", X"1D60",            "----------------", X"1D64",            "----------------",
		X"1D68",            "----------------", X"1D6C",            "----------------", X"1D71",
		"----------------", X"1D75",            X"1D76",            "----------------", X"1D77",
		X"1D78",            "----------------", X"1D79",            X"1D7A",            X"1D7B",            X"1D7C", -- CPSE bubble inserted
		X"1D7D",            "----------------", "----------------", "----------------", X"1D7E",            "----------------", X"1D84",            "----------------", -- ADD bubble inserted (x3)
		X"1D88",            "----------------", X"1D8B",            "----------------", X"1D9F",
		"----------------", X"1DA4",            "----------------", X"1DA8",            X"1DA9",
		"----------------", X"1DAA",            X"1DAB",            "----------------", X"1DAC",            X"1DAD", -- CPSE bubble inserted
		X"1DAE",            X"1DAF",            "----------------", "----------------", "----------------", X"1DB0",            "----------------", X"1DB2", -- ADD bubble inserted (x3)
		"----------------", X"1DB6",            "----------------", X"1DBA",            "----------------",
		X"1DBF",            "----------------", X"1DC4",            "----------------", X"1DC8",
		X"1DC9",            "----------------", X"1DCA",            X"1DCB",            "----------------", X"1DCC", -- CPSE bubble inserted
		X"1DCD",            X"1DCE",            X"1DCF",            "----------------", "----------------", "----------------", X"1DD0",            "----------------", -- ADD bubble inserted (x3)
		X"1DD2",            "----------------", X"1DD6",            "----------------", X"1DDA",
		"----------------", X"1DDE",            "----------------", X"1DE2",            "----------------",
		X"1DE6",            X"1DE7",            "----------------", X"1DE8",            X"1DE9",            "----------------", -- CPSE bubble inserted
		X"1DEA",            X"1DEB",            X"1DEC",            X"1DED",            X"1DEE",            "----------------", "----------------", "----------------", -- ADIW bubble inserted (x3)
		"----------------", X"1DEF",            "----------------", X"1DF4",            "----------------",
		X"1DF8",            "----------------", X"1DFB",            "----------------", X"1DFF",
		"----------------", X"1E04",            X"1E05",            "----------------", X"1E06",
		X"1E07",            "----------------", X"1E08",            X"1E09",            X"1E0A",            "----------------", -- CPSE bubble inserted
		X"1E0B",            X"1E0C",            X"1E0D",            "----------------", X"1E0E",            X"1E0F", -- CPSE bubble inserted
		X"1E10",            X"1E11",            X"1E12",            "----------------", "----------------", "----------------", "----------------", X"1E13", -- ADIW bubble inserted (x3)
		"----------------", X"1E16",            "----------------", X"1E1A",            "----------------",
		X"1E1E",            "----------------", X"1E23",            "----------------", X"1E27",
		X"1E28",            "----------------", X"1E29",            X"1E2A",            "----------------",
		X"1E2B",            X"1E2C",            X"1E2D",            "----------------", X"1E2E",            X"1E2F", -- CPSE bubble inserted
		X"1E30",            "----------------", X"1E31",            X"1E32",            X"1E33",            X"1E34", -- CPSE bubble inserted
		X"1E35",            "----------------", "----------------", "----------------", "----------------", X"1E36",            "----------------", X"1E40", -- ADIW bubble inserted (x3)
		"----------------", X"1E44",            "----------------", X"1E48",            "----------------",
		X"1E4B",            "----------------", X"1E4F",            X"1E50",            "----------------",
		X"1E51",            X"1E52",            "----------------", X"1E53",            X"1E54",
		X"1E55",            "----------------", X"1E56",            X"1E57",            X"1E58",            "----------------", X"1E59", -- CPSE bubble inserted (x2)
		X"1E5A",            X"1E5B",            X"1E5C",            X"1E5D",            "----------------", "----------------", "----------------", X"1E5E", -- AND bubble inserted (x3)
		"----------------", X"1E62",            "----------------", X"1E66",            "----------------",
		X"1E6A",            "----------------", X"1E6F",            X"1E70",            "----------------",
		X"1E71",            X"1E72",            "----------------", X"1E73",            X"1E74",            X"1E75", -- CPSE bubble inserted
		X"1E76",            "----------------", "----------------", "----------------", X"1E77",            "----------------", X"1E7A",            "----------------", -- AND bubble inserted (x3)
		X"1E7F",            "----------------", X"1E84",            "----------------", X"1E88",
		X"1E89",            "----------------", X"1E8A",            X"1E8B",            "----------------", X"1E8C", -- CPSE bubble inserted
		X"1E8D",            X"1E8E",            X"1E8F",            "----------------", "----------------", "----------------", X"1E90",            "----------------", -- AND bubble inserted (x3)
		X"1E94",            "----------------", X"1E98",            "----------------", X"1E9B",
		"----------------", X"1E9F",            X"1EA0",            "----------------", X"1EA1",
		X"1EA2",            "----------------", X"1EA3",            X"1EA4",            X"1EA5",            X"1EA6", -- CPSE bubble inserted
		"----------------", "----------------", "----------------", X"1EA7",            "----------------", X"1EAD",            "----------------", X"1EB2", -- ANDI bubble inserted (x3)
		"----------------", X"1EB6",            "----------------", X"1EBB",            X"1EBC",
		"----------------", X"1EBD",            X"1EBE",            "----------------", X"1EBF",            X"1EC0", -- CPSE bubble inserted
		X"1EC1",            "----------------", "----------------", "----------------", X"1EC2",            "----------------", X"1EC8",            "----------------", -- ANDI bubble inserted (x3)
		X"1ECB",            "----------------", X"1ECF",            "----------------", X"1ED4",
		X"1ED5",            "----------------", X"1ED6",            X"1ED7",            "----------------", X"1ED8", -- CPSE bubble inserted
		X"1ED9",            X"1EDA",            "----------------", "----------------", "----------------", X"1EDB",            "----------------", X"1EDF", -- ANDI bubble inserted (x3)
		"----------------", X"1EE2",            "----------------", X"1EE6",            "----------------",
		X"1EEB",            X"1EEC",            "----------------", X"1EED",            X"1EEE",            "----------------", -- CPSE bubble inserted
		X"1EEF",            X"1EF0",            X"1EF1",            X"1EF2",            "----------------", "----------------", "----------------", X"1EF3", -- ASR bubble inserted (x3)
		"----------------", X"1EF6",            "----------------", X"1EFB",            "----------------",
		X"1EFF",            "----------------", X"1F03",            "----------------", X"1F06",
		X"1F07",            "----------------", X"1F08",            X"1F09",            "----------------", X"1F0A", -- CPSE bubble inserted
		X"1F0B",            X"1F0C",            X"1F0D",            "----------------", "----------------", "----------------", X"1F0E",            "----------------", -- ASR bubble inserted (x3)
		X"1F14",            "----------------", X"1F18",            "----------------", X"1F1B",
		"----------------", X"1F1E",            "----------------", X"1F22",            X"1F23",
		"----------------", X"1F24",            X"1F25",            "----------------", X"1F26",            X"1F27", -- CPSE bubble inserted
		X"1F28",            X"1F29",            "----------------", "----------------", "----------------", X"1F2A",            "----------------", X"1F2D", -- ASR bubble inserted (x3)
		"----------------", X"1F32",            "----------------", X"1F36",            "----------------",
		X"1F3B",            "----------------", X"1F3F",            X"1F40",            "----------------",
		X"1F41",            X"1F42",            "----------------", X"1F43",            X"1F44",            X"1F45", -- CPSE bubble inserted
		"----------------", "----------------", "----------------", X"1F46",            "----------------", X"1F4A",            "----------------", "----------------", "----------------", X"1F4B",            "----------------", 
		X"1F4E",            "----------------", "----------------", "----------------", X"1F4F",            "----------------", X"1F52",            "----------------", "----------------", "----------------", X"1F53",
		"----------------", X"1F56",            "----------------", "----------------", "----------------", X"1F57",            "----------------", X"1F5B", "----------------", "----------------", "----------------", 
		X"1F5C",            "----------------", X"1F5F",            "----------------", "----------------", "----------------", X"1F60",            "----------------",
		X"1F64",            "----------------", "----------------", "----------------", X"1F65",            "----------------", X"1F68",            "----------------", "----------------", "----------------", X"1F69",
		"----------------", X"1F6C",            "----------------", "----------------", "----------------", X"1F6D",            "----------------", X"1F72", "----------------", "----------------", "----------------", 
		X"1F73",            "----------------", X"1F76",            "----------------", "----------------", "----------------", X"1F77",            "----------------",
		X"1F7B",            "----------------", "----------------", "----------------", X"1F7C",            "----------------", X"1F7F",            "----------------", "----------------", "----------------", X"1F80",
		"----------------", X"1F83",            "----------------", "----------------", "----------------", X"1F84",            "----------------", X"1F87",
		"----------------", "----------------", "----------------", X"1F88",            "----------------", X"1F8C",            X"1F8D",            X"1F8E", "----------------", "----------------", "----------------", 
		X"1F8F",            "----------------", X"1F93",            "----------------", "----------------", "----------------", X"1F94",            X"1F95", "----------------", 
		X"1F96",            X"1F97",            X"1F98",            "----------------", "----------------", "----------------", X"1F99",            "----------------",
		X"1F9D",            "----------------", "----------------", "----------------", X"1F9E",            X"1F9F",            "----------------", X"1FA0",            X"1FA1",
		X"1FA2",            X"1FA3",            "----------------", "----------------", "----------------", X"1FA4",            "----------------", X"1FA8",
		"----------------", X"1FAC",            "----------------", X"1FB0",            "----------------",
		X"1FB4",            "----------------", X"1FB8",            X"1FB9",            "----------------",
		X"1FBA",            X"1FBB",            "----------------", X"1FBC",            X"1FBD",            X"1FBE",
		X"1FBF",            "----------------", "----------------", "----------------", X"1FC0",            "----------------", X"1FC2",            "----------------",
		X"1FC6",            "----------------", X"1FCA",            "----------------", X"1FCE",
		"----------------", X"1FD2",            X"1FD3",            "----------------", X"1FD4",
		X"1FD5",            "----------------", X"1FD6",            X"1FD7",            X"1FD8",            X"1FD9", "----------------", "----------------", "----------------", 
		X"1FDA",            "----------------", X"1FDD",            "----------------", X"1FE2",
		"----------------", X"1FE6",            "----------------", X"1FEA",            "----------------",
		X"1FEE",            X"1FEF",            "----------------", X"1FF0",            X"1FF1", "----------------", 
		X"1FF2",            X"1FF3",            X"1FF4",            X"1FF5",            X"1FF6", "----------------", "----------------", "----------------", 
		X"1FF7",            "----------------", X"1FFB",            "----------------", X"1FFF",
		"----------------", X"2004",            "----------------", X"2008",            "----------------",
		X"200B",            "----------------", X"200E",            X"200F",            "----------------",
		X"2010",            X"2011",            X"2012",            "----------------", "----------------", "----------------", X"2013",            "----------------",
		X"2018",            "----------------", X"201B",            "----------------", X"201E",
		"----------------", X"2022",            "----------------", X"2026",            "----------------",
		X"202A",            X"202B",            "----------------", X"202C",            X"202D",
		X"202E",            "----------------", "----------------", "----------------", X"202F",            "----------------", X"2034",            "----------------",
		X"2038",            "----------------", X"203B",            "----------------", X"203F",
		"----------------", X"2042",            "----------------", X"2046",            X"2047",
		"----------------", X"2048",            X"2049",            X"204A",            "----------------", "----------------", "----------------", X"204B", "----------------", "----------------", "----------------", 
		X"204C",            "----------------", X"2050",            "----------------", X"2054",
		"----------------", X"2058",            "----------------", X"205B",            "----------------",
		X"205E",            "----------------", X"2062",            X"2063",            "----------------",
		X"2064",            X"2065",            X"2066",            "----------------", "----------------", "----------------", X"2067",            "----------------", "----------------", "----------------", X"2068",
		"----------------", X"206C",            "----------------", X"206F",            "----------------",
		X"2074",            "----------------", X"2078",            "----------------", X"207B",
		"----------------", X"207E",            X"207F",            "----------------", X"2080",
		X"2081",            X"2082",            "----------------", "----------------", "----------------", X"2083",            "----------------", "----------------", "----------------", X"2084",            "----------------", "----------------", "----------------", X"2085",
		"----------------", X"208A",            "----------------", X"208E",            "----------------",
		X"2092",            "----------------", X"2096",            "----------------", X"209A",
		"----------------", X"209E",            X"209F",            "----------------", X"20A0",
		X"20A1",            "----------------", "----------------", "----------------", X"20A2",            "----------------", X"20A6",            "----------------",
		X"20AA",            "----------------", X"20AE",            "----------------", X"20B2",
		"----------------", X"20B6",            "----------------", X"20BA",            X"20BB",
		"----------------", X"20BC",            X"20BD",            "----------------", "----------------", "----------------", X"20BE",            "----------------",
		X"20C2",            "----------------", X"20C6",            "----------------", X"20CA",
		"----------------", X"20CE",            "----------------", X"20D2",            "----------------",
		X"20D6",            X"20D7",            "----------------", X"20D8",            X"20D9",            "----------------", "----------------", "----------------", 
		X"20DA",            "----------------", X"20E0",            "----------------", X"20E4",
		"----------------", X"20E8",            "----------------", X"20EB",            "----------------",
		X"20EF",            "----------------", X"20F3",            X"20F4",            "----------------",
		X"20F5",            X"20F6",            "----------------", "----------------", "----------------", X"20F7",            "----------------", X"20FB",
		"----------------", X"20FF",            "----------------", X"2104",            "----------------",
		X"2108",            X"2109",            "----------------", X"210A",            X"210B",            "----------------", 
		X"210C",            X"210D",            X"210E",            "----------------", "----------------", "----------------", X"210F",            "----------------", "----------------", "----------------", X"2110",
		"----------------", X"2114",            "----------------", X"2118",            "----------------",
		X"211C",            "----------------", X"211F",            X"2120",            "----------------",
		X"2121",            X"2122",            "----------------", X"2123",            X"2124",            X"2125",
		X"2126",            X"2127",            "----------------", "----------------", "----------------", X"2128",            "----------------", X"212B",
		"----------------", X"212F",            "----------------", X"2134",            "----------------",
		X"2138",            X"2139",            "----------------", X"213A",            X"213B",            "----------------", 
		X"213C",            X"213D",            X"213E",            X"213F",            X"2140",            "----------------", "----------------", "----------------", 
		X"2141",            "----------------", X"2144",            "----------------", X"2148",
		"----------------", X"214B",            "----------------", X"214F",            X"2150",
		"----------------", X"2151",            X"2152",            "----------------", X"2153",            X"2154",
		X"2155",            X"2156",            X"2157",            "----------------", "----------------", "----------------", X"2158",            "----------------",
		X"215C",            "----------------", X"215F",            "----------------", X"2164",
		"----------------", X"2168",            X"2169",            "----------------", X"216A",
		X"216B",            "----------------", X"216C",            X"216D",            X"216E",            X"216F", "----------------", "----------------", "----------------", 
		X"2170",            "----------------", X"2174",            "----------------", X"2178",
		"----------------", X"217B",            "----------------", X"217F",            "----------------",
		X"2184",            X"2185",            "----------------", X"2186",            X"2187", "----------------", 
		X"2188",            X"2189",            X"218A",            X"218B",            "----------------", "----------------", "----------------", X"218C",
		"----------------", X"218F",            "----------------", X"2194",            "----------------",
		X"2198",            "----------------", X"219B",            "----------------", X"219F",
		X"21A0",            "----------------", X"21A1",            X"21A2",            "----------------", X"21A3",
		X"21A4",            X"21A5",            X"21A6",            "----------------", "----------------", "----------------", X"21A7",            "----------------",
		X"21AA",            "----------------", X"21AE",            "----------------", X"21B4",
		"----------------", X"21B8",            "----------------", X"21BB",            X"21BC",
		"----------------", X"21BD",            X"21BE",            "----------------", X"21BF",            X"21C0",
		X"21C1",            X"21C2",            "----------------", "----------------", "----------------", X"21C3",            "----------------", X"21C8",
		"----------------", X"21CB",            "----------------", X"21CF",            "----------------",
		X"21D4",            "----------------", X"21D8",            X"21D9",            "----------------",
		X"21DA",            X"21DB",            "----------------", X"21DC",            X"21DD",            X"21DE",
		X"21DF",            "----------------", "----------------", "----------------", X"21E0",            "----------------", X"21E4",            "----------------",
		X"21E8",            "----------------", X"21EB",            "----------------", X"21EF",
		"----------------", X"21F4",            X"21F5",            "----------------", X"21F6",
		X"21F7",            "----------------", X"21F8",            X"21F9",            X"21FA",            X"21FB", "----------------", "----------------", "----------------", 
		X"21FC",            "----------------", X"2202",            "----------------", X"2206",
		"----------------", X"220A",            "----------------", X"220E",            "----------------",
		X"2214",            X"2215",            "----------------", X"2216",            X"2217", "----------------", 
		X"2218",            X"2219",            X"221A",            X"221B",            X"221C", "----------------", "----------------", "----------------", 
		X"221D",            "----------------", X"2224",            "----------------", X"2228",
		"----------------", X"222B",            "----------------", X"222F",            X"2230",
		"----------------", X"2231",            X"2232",            "----------------", X"2233",            X"2234",
		X"2235",            X"2236",            X"2237",            "----------------", "----------------", "----------------", X"2238",            "----------------",
		X"223D",            "----------------", X"2242",            "----------------", X"2246",
		"----------------", X"224A",            X"224B",            "----------------", X"224C",
		X"224D",            "----------------", X"224E",            X"224F",            X"2250",            X"2251",
		X"2252",            "----------------", "----------------", "----------------", X"2253",            "----------------", X"2258",            "----------------",
		X"225B",            "----------------", X"225E",            "----------------", X"2262",
		X"2263",            "----------------", X"2264",            X"2265",            "----------------", X"2266",
		X"2267",            X"2268",            X"2269",            "----------------", "----------------", "----------------", X"226A",            "----------------",
		X"226E",            "----------------", X"2272",            "----------------", X"2276",
		"----------------", X"227A",            X"227B",            "----------------", X"227C",
		X"227D",            "----------------", X"227E",            X"227F",            X"2280",            X"2281", "----------------", "----------------", "----------------", 
		X"2282",            "----------------", X"2286",            "----------------", X"228A",
		"----------------", X"228E",            "----------------", X"2292",            X"2293",
		"----------------", X"2294",            X"2295",            "----------------", X"2296",            X"2297",
		X"2298",            X"2299",            "----------------", "----------------", "----------------", X"229A",            "----------------", X"229F",
		"----------------", X"22A4",            "----------------", X"22A8",            "----------------",
		X"22AB",            X"22AC",            "----------------", X"22AD",            X"22AE", "----------------", 
		X"22AF",            X"22B0",            X"22B1",            "----------------", "----------------", "----------------", X"22B2",            X"22B3", "----------------", "----------------", "----------------", 
		X"22B4",            "----------------", X"22B8",            "----------------", X"22BB",
		"----------------", X"22BE",            "----------------", X"22C4",            "----------------",
		X"22C8",            X"22C9",            "----------------", X"22CA",            X"22CB", "----------------", 
		X"22CC",            X"22CD",            X"22CE",            X"22CF",            "----------------", "----------------", "----------------", X"22D0",
		"----------------", X"22D4",            "----------------", X"22D8",            "----------------",
		X"22DB",            "----------------", X"22DE",            "----------------", X"22E2",
		X"22E3",            "----------------", X"22E4",            X"22E5",            "----------------", X"22E6",
		X"22E7",            X"22E8",            X"22E9",            "----------------", "----------------", "----------------", X"22EA",            "----------------",
		X"22EE",            "----------------", X"22F2",            "----------------", X"22F6",
		"----------------", X"22FA",            "----------------", X"22FE",            X"22FF",
		"----------------", X"2300",            X"2301",            "----------------", X"2302",            X"2303",
		X"2304",            "----------------", "----------------", "----------------", X"2305",            X"2306",            X"2307",            "----------------", "----------------", "----------------", X"2308",
		"----------------", X"230E",            "----------------", X"2312",            "----------------",
		X"2316",            "----------------", X"231A",            "----------------", X"231E",
		"----------------", X"2322",            X"2323",            "----------------", X"2324",
		X"2325",            "----------------", X"2326",            X"2327",            X"2328",            X"2329", "----------------", "----------------", "----------------", 
		X"232A",            "----------------", X"232E",            "----------------", X"2332",
		"----------------", X"2336",            "----------------", X"233A",            "----------------",
		X"233E",            "----------------", X"2342",            X"2343",            "----------------",
		X"2344",            X"2345",            "----------------", X"2346",            X"2347",            X"2348",
		X"2349",            "----------------", "----------------", "----------------", X"234A",            "----------------", X"234E",            "----------------",
		X"2352",            "----------------", X"2356",            "----------------", X"235A",
		"----------------", X"235E",            "----------------", X"2362",            X"2363",
		"----------------", X"2364",            X"2365",            "----------------", X"2366",            X"2367",
		X"2368",            "----------------", "----------------", "----------------", X"2369",            X"236A",            "----------------", "----------------", "----------------", X"236B",            "----------------",
		X"2372",            "----------------", X"2376",            "----------------", X"237A",
		"----------------", X"237E",            "----------------", X"2382",            "----------------",
		X"2386",            X"2387",            "----------------", X"2388",            X"2389", "----------------", 
		X"238A",            X"238B",            X"238C",            X"238D",            "----------------", "----------------", "----------------", X"238E",
		"----------------", X"2394",            "----------------", X"2398",            "----------------",
		X"239B",            "----------------", X"239E",            "----------------", X"23A2",
		"----------------", X"23A6",            X"23A7",            "----------------", X"23A8",
		X"23A9",            "----------------", X"23AA",            X"23AB",            X"23AC",            X"23AD", "----------------", "----------------", "----------------", 
		X"23AE",            "----------------", X"23B4",            "----------------", X"23B8",
		"----------------", X"23BB",            "----------------", X"23BE",            "----------------",
		X"23C2",            "----------------", X"23C6",            X"23C7",            "----------------",
		X"23C8",            X"23C9",            "----------------", X"23CA",            X"23CB",            X"23CC",
		X"23CD",            X"23CE",            "----------------", "----------------", "----------------", "----------------", X"23CF",            "----------------",
		X"23D4",            "----------------", X"23D8",            "----------------", X"23DB",
		"----------------", X"23DE",            "----------------", X"23E2",            X"23E3",
		"----------------", X"23E4",            X"23E5",            "----------------", X"23E6",
		X"23E7",            X"23E8",            "----------------", X"23E9",            X"23EA",            X"23EB", "----------------", 
		X"23EC",            X"23ED",            X"23EE",            X"23EF",            X"23F0", "----------------", "----------------", "----------------", 
		"----------------", X"23F1",            "----------------", X"23F6",            "----------------",
		X"23FA",            "----------------", X"23FE",            "----------------", X"2402",
		"----------------", X"2406",            X"2407",            "----------------", X"2408",
		X"2409",            "----------------", X"240A",            X"240B",            X"240C", "----------------", 
		X"240D",            X"240E",            X"240F",            "----------------", X"2410",            X"2411",
		X"2412",            X"2413",            X"2414",            "----------------", "----------------", "----------------", "----------------", X"2415",
		"----------------", X"241A",            "----------------", X"241E",            "----------------",
		X"2422",            "----------------", X"2426",            "----------------", X"242A",
		X"242B",            "----------------", X"242C",            X"242D",            "----------------",
		X"242E",            X"242F",            X"2430",            "----------------", X"2431",            X"2432",
		X"2433",            "----------------", X"2434",            X"2435",            X"2436",            X"2437",
		X"2438",            "----------------", "----------------", "----------------", X"2439",            "----------------", X"243E",            "----------------",
		X"2442",            "----------------", X"2446",            "----------------", X"244A",
		"----------------", X"244E",            "----------------", X"2452",            X"2453",
		"----------------", X"2454",            X"2455",            "----------------", X"2456",            X"2457",
		X"2458",            X"2459",            "----------------", "----------------", "----------------", X"245A",            "----------------", X"245E",
		"----------------", X"2462",            "----------------", X"2466",            "----------------",
		X"247A",            "----------------", X"247E",            "----------------", X"2482",
		X"2483",            "----------------", X"2484",            X"2485",            "----------------", X"2486",
		X"2487",            X"2488",            X"2489",            "----------------", "----------------", "----------------", X"248A",            "----------------",
		X"248E",            "----------------", X"2492",            "----------------", X"2496",
		"----------------", X"249A",            "----------------", X"249E",            "----------------",
		X"24A2",            X"24A3",            "----------------", X"24A4",            X"24A5", "----------------", 
		X"24A6",            X"24A7",            X"24A8",            X"24A9",            "----------------", "----------------", "----------------", X"24AA",
		"----------------", X"24AE",            "----------------", X"24B2",            "----------------",
		X"24B6",            "----------------", X"24BA",            "----------------", X"24BE",
		"----------------", X"24C2",            X"24C3",            "----------------", X"24C4",
		X"24C5",            "----------------", X"24C6",            X"24C7",            X"24C8",            X"24C9", "----------------", "----------------", "----------------", 
		X"24CA",            "----------------", X"24CE",            "----------------", X"24D2",
		"----------------", X"24D6",            "----------------", X"24DA",            "----------------",
		X"24DE",            "----------------", X"24E2",            X"24E3",            "----------------",
		X"24E4",            X"24E5",            "----------------", X"24E6",            X"24E7",            X"24E8",
		X"24E9",            "----------------", "----------------", "----------------", X"24EA",            "----------------", X"24EE",            "----------------",
		X"24F2",            "----------------", X"24F6",            "----------------", X"24FA",
		"----------------", X"24FE",            "----------------", X"2502",            X"2503",
		"----------------", X"2504",            X"2505",            "----------------", X"2506",            X"2507",
		X"2508",            X"2509",            X"250A",            X"250B",            "----------------", X"250C",
		X"250D",            X"250E",            X"250F",            X"2510",            X"2511", "----------------", 
		X"2512",            X"2513",            X"2514",            X"2515",            X"2516",
		X"2517",            "----------------", X"2518",            X"2519",            X"251A",            X"251B",
		X"251C",            "----------------", "----------------", "----------------", "----------------", X"251D",            "----------------", X"2540",
		"----------------", X"2544",            X"2545",            X"2546",            "----------------", X"2547",
		X"2548",            X"2549",            "----------------", X"254A",            X"254B",            X"254C",
		X"254D",            X"254E",            "----------------", "----------------", "----------------", "----------------", X"254F",            "----------------",
		X"2560",            "----------------", X"2564",            X"2565",            X"2566", "----------------", 
		X"2567",            X"2568",            X"2569",            "----------------", X"256A",            X"256B",
		X"256C",            X"256D",            X"256E",            "----------------", "----------------", "----------------", "----------------", X"256F",
		"----------------", X"2580",            "----------------", X"2584",            X"2585",
		X"2586",            "----------------", X"2587",            X"2588",            X"2589",            "----------------", X"258A",
		X"258B"
		);

	-- Data Read Vector
	constant DataReadTest : std_logic_vector(0 to 2764) := 
		"11111111111111111111111101111111110111111111011111111101111111111111111111111111111111111111111111111111111110111111110111111101111111111111111111111111111101111111101111111101111111111111111111111111111101111111101111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111001111111111110011111111111100111111111111110011111111111111001111111111111111001111111111111111100111111111111111101111111111011111111110111111111101111111111011111111110111111111101111111111011111111110111111111101111111111011111111110111111111101111111111011111111110111111111101111111110111111111011111111101111111110111111111011111111101111111110111111111011111111101111111110111111111011111111101111111110111111111011111111101111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";

	-- Data Write Vector
	constant DataWriteTest : std_logic_vector(0 to 2764) := 
		"11111011101110111011101111101110111110111011111011101111101111011110111101111011111101111101111101111101111011101110111101110111011111101110111110111011110111011101111011101111011111101110111110111011110111011101111011101111011111101110111110111011111011101111101110111110111011111011101111101110111110111011111011101111101110111110111011111011101101110111110101011111110110110111110111111111011111111101111111111111011111111101111111110111111111110111111111111101111110111111011111011111011111110111111101110011011111101110011011111101100110111111011001101111110111100110111111011110011011111101111111110011111111101111111001111111110111111101111111111011111111110111111111101111111111011111111110111111111101111111111011111111110111111111101111111111011111111110111111111101111111111011111111110111111111101111111110111111111011111111101111111110111111111011111111101111111110111111111011111111101111111110111111111011111111101111111110111111111011111111101111111110111111111111111111111111111101111111111111111111111110111111111111111111111111011111111111111111111111110111111111111111111111111011111111111111111111111101111111111111111111111110110111111111111111111111111111110110111111111111111111111111111110110111111111111111111111111110111111111111111111110111111111111111111110111111111111111111110111111111111111111101111111111111111111011111111111111111111110111111111111111111111101111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111011111111111111111111110111111111111111111111111101111111111111111111101111111111111111111101111111111111111111111110111111111111111111111111011111111111111111111111111110111111111111111111101111111111111111111011111111111111111110111111111111111011111111111111111111111011111111111111111111101111111111111111111110111111111111111111111011111111111111111111110111111111111111111111101111111111111111111111011111111111111111111110111111111111111111111101111111111111111111111011111111111111111111101111111111111111111110111111111111111111111011111111111111111111011111111111111111111011111111111111111111011111111111111111111111111011111111111111111111110111111111111111111111101111111111111111111111111111101111111111111111111111110111111111111111111111111011111111111111111111111111110111111111111111111111111011111111111111111111111101111111111111111111111110110111111111111111111111111111110110111111111111111111111111111110110111111111111111111111111111111011111111111111111111111101111111111111111111111110111111111111111111111111011111111111111111111111101111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";

	-- Data Data Bus Test In Vectors
	constant DataDBTestIn : testarray2 := (
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", X"45",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", X"F0",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", X"11",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", X"00",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", X"21",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		X"4A",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"00",      "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"21",      "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", X"4A",      "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", X"00",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", X"21",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		X"2B",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"03",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", X"67",      "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", X"8F",      "ZZZZZZZZ", X"A5",      "ZZZZZZZZ",
		X"80",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", -- SBRS/SBRC bubbles
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", -- CPSE bubbles
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		X"E1",      X"14",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		X"E6",      X"14",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"EA",
		X"14",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"EE",      X"14",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"F4",
		X"14",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		X"FA",      X"14",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		X"24",      X"1A",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", X"39",      X"1A",      "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"FF",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"01",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"02",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"03",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"04",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"05",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"06",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"07",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"08",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"09",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"10",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"11",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"12",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"13",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"14",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"15",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"16",      "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", X"17",      "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", X"18",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		X"19",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"20",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"21",      "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", X"22",      "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", X"23",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		X"24",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"25",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"26",      "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", X"27",      "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", X"28",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		X"29",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"30",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"31",      "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",  "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ",
		"ZZZZZZZZ"
	);

	-- Data Data Bus Test Out Vectors
	constant DataDBTestOut : testarray2 := (
		"--------", "--------", "--------", "--------", "--------", X"23",      "--------", "--------",
		"--------", X"FF",      "--------", "--------", "--------",
		X"01",      "--------", "--------", "--------", X"00",
		"--------", "--------", "--------", X"45",      "--------",
		"--------", "--------", "--------", "--------", X"45",
		"--------", "--------", "--------", X"F0",      "--------",
		"--------", "--------", "--------", "--------", X"F0",
		"--------", "--------", "--------", X"11",      "--------",
		"--------", "--------", "--------", "--------", X"11",
		"--------", "--------", "--------", X"00",      "--------",
		"--------", "--------", "--------", "--------", X"00",
		"--------", "--------", "--------", "--------", X"CD",
		"--------", "--------", "--------", "--------", X"90",
		"--------", "--------", "--------", "--------", X"13",
		"--------", "--------", "--------", "--------", X"00",
		"--------", "--------", "--------", "--------", "--------",
		"--------", X"89",      "--------", "--------", "--------",
		"--------", "--------", X"44",      "--------", "--------",
		"--------", "--------", "--------", X"89",      "--------",
		"--------", "--------", "--------", "--------", X"00",
		"--------", "--------", "--------", "--------", X"21",
		"--------", "--------", "--------", X"21",      "--------",
		"--------", "--------", X"4A",      "--------", "--------",
		"--------", "--------", X"4A",      "--------", "--------",
		"--------", X"00",      "--------", "--------", "--------",
		X"00",      "--------", "--------", "--------", "--------",
		"--------", "--------", X"32",      "--------", "--------",
		"--------", X"DA",      "--------", "--------", "--------",
		"--------", "--------", X"56",      "--------", "--------",
		"--------", X"07",      "--------", "--------", "--------",
		"--------", X"21",      "--------", "--------", "--------",
		X"21",      "--------", "--------", "--------", X"4A",
		"--------", "--------", "--------", "--------", X"4A",
		"--------", "--------", "--------", X"00",      "--------",
		"--------", "--------", "--------", X"00",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		X"01",      "--------", "--------", "--------", X"43",
		"--------", "--------", "--------", "--------", "--------",
		X"1F",      "--------", "--------", "--------", X"76",
		"--------", "--------", "--------", "--------", X"21",
		"--------", "--------", "--------", X"21",      "--------",
		"--------", "--------", X"2B",      "--------", "--------",
		"--------", "--------", X"2B",      "--------", "--------",
		"--------", X"03",      "--------", "--------", "--------",
		"--------", X"03",      "--------", "--------", "--------",
		"--------", "--------", "--------", X"32",      "--------",
		"--------", "--------", X"DA",      "--------", "--------",
		"--------", "--------", "--------", X"56",      "--------",
		"--------", "--------", X"07",      "--------", "--------",
		"--------", "--------", "--------", X"01",      "--------",
		"--------", "--------", X"43",      "--------", "--------",
		"--------", "--------", "--------", X"1F",      "--------",
		"--------", "--------", X"76",      "--------", "--------",
		"--------", "--------", "--------", X"4D",      "--------",
		"--------", "--------", X"EA",      "--------", "--------",
		"--------", "--------", "--------", X"3E",      "--------",
		"--------", "--------", X"6B",      "--------", "--------",
		"--------", "--------", "--------", X"32",      "--------",
		"--------", "--------", X"DA",      "--------", "--------",
		"--------", "--------", "--------", X"56",      "--------",
		"--------", "--------", X"07",      "--------", "--------",
		"--------", "--------", "--------", X"01",      "--------",
		"--------", "--------", X"43",      "--------", "--------",
		"--------", "--------", "--------", X"1F",      "--------",
		"--------", "--------", X"76",      "--------", "--------",
		"--------", "--------", "--------", X"4D",      "--------",
		"--------", "--------", X"EA",      "--------", "--------",
		"--------", "--------", "--------", X"3E",      "--------",
		"--------", "--------", X"6B",      "--------", "--------",
		X"67",      "--------", "--------", "--------", X"67",
		"--------", "--------", "--------", "--------", "--------",
		X"80",      "--------", X"A5",      "--------", X"8F",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"8F",      "--------", "--------",
		X"A5",      "--------", "--------", X"80",      "--------",
		"--------", "--------", "--------", "--------", X"A5",      "--------", "--------", -- SBRC bubbles (x2)
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"04",      "--------", "--------", "--------", "--------", -- SBRC bubbles (x2)
		"--------", "--------", "--------", "--------", "--------", X"95",      "--------", -- SBRC bubbles (x2)
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", -- SBRS bubbles (x2)
		X"66",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", X"BE",      "--------", -- SBRS bubbles (x2)
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"01",      "--------", "--------", "--------", -- SBRS bubbles (x2)
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", -- CPSE bubbles (x2)
		"--------", X"FF",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", -- CPSE bubbles (x3)
		"--------", "--------", X"37",      "--------", "--------",
		"--------", "--------", "--------", "--------", X"55",
		"--------", "--------", "--------", "--------", "--------",
		"--------", X"2C",      "--------", "--------", "--------",
		"--------", "--------", X"44",      "--------", "--------",
		"--------", "--------", "--------", X"01",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", X"99",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"20",
		"--------", "--------", "--------", X"14",      "--------",
		"--------", "--------", X"8E",      "--------", "--------",
		"--------", "--------", "--------", "--------", X"8E",
		"--------", "--------", "--------", X"14",      "--------",
		"--------", "--------", X"22",      "--------", "--------",
		"--------", "--------", "--------", "--------", X"22",
		"--------", "--------", X"14",      X"EA",      "--------",
		"--------", X"45",      "--------", "--------", "--------",
		"--------", "--------", "--------", X"45",      "--------",
		"--------", X"14",      X"EE",      "--------", "--------",
		X"EA",      "--------", "--------", "--------", "--------",
		"--------", "--------", X"EA",      "--------", "--------",
		"--------", "--------", X"14",      X"F4",      "--------", 
		"--------", X"07",      "--------", "--------", "--------",
		"--------", "--------", "--------", X"07",      "--------",
		"--------", "--------", "--------", X"14",      X"FA",
		"--------", "--------", X"11",      "--------", "--------",
		"--------", "--------", "--------", "--------", X"11",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"1A",      X"24",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"99",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"1A",      X"39",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"E0",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", X"FF",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"01",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"02",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"03",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"04",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"05",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"06",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"07",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"08",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"09",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"10",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"11",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"12",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"13",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"14",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"15",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		X"16",      "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", X"17",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", X"18",      "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", X"19",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"20",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		X"21",      "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", X"22",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", X"23",      "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", X"24",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"25",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		X"26",      "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", X"27",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", X"28",      "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", X"29",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"30",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		X"31",      "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		X"9A",      "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"2C",      "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", X"D3",      "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", X"9A",
		"--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		X"2C",      "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", X"D2",      "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", X"7F",      "--------", "--------",
		X"5A",      "--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		X"01",      "--------", "--------", X"00",      "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", X"3D",      "--------",
		"--------", X"00",      "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"40",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		X"52",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"00",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"4D",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		X"00",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"00",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		X"DB",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"2C",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"FF",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", 
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"8C",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"FF",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"AA",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"73",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"04",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"55",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"73",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"04",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"04",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"40",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", X"08",      "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"91",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"FE",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"00",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"9F",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"B1",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"87",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"7B",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		X"2A",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"3C",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"0A",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"AB",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"88",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"F6",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"7F",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		X"FF",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"FF",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"57",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"78",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"7B",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		X"2A",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"BC",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"E6",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"77",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"1E",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"DA",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"AE",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"79",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"01",
		"--------", "--------", X"5A",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"FD",      "--------", "--------",
		X"FF",      "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		X"C1",      "--------", "--------", X"FF",      "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"E6",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		X"78",      "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", X"1E",      "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", X"41",      "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", X"5B",      "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", X"78",      "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------", "--------", "--------", "--------", "--------",
		"--------"
	);


	-- Data Address Bus Test Vectors
	constant DataABTest : testarray := (
		"----------------", "----------------", "----------------", "----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------",
		X"1000",            "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", X"1000",            "----------------", "----------------", X"0900",
		"----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", X"1000",            "----------------", "----------------", X"0900",
		"----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", X"1000",            "----------------", "----------------", X"0900",
		"----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", X"1000",            "----------------", "----------------", X"0900",
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"BBAA",            "----------------", "----------------", "----------------",
		"----------------", "----------------", X"FA01",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"FFFF",            "----------------",
		"----------------", "----------------", "----------------", "----------------", X"0001",
		"----------------", "----------------", "----------------", "----------------", X"0FFF",
		"----------------", X"0FFF",            "----------------", X"0900",            "----------------",
		"----------------", "----------------", X"0FFF",            "----------------", "----------------",
		X"0FFF",            "----------------", X"0900",            "----------------", "----------------",
		"----------------", X"0FFF",            "----------------", X"0FFF",            "----------------",
		X"0900",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"11A0",            "----------------", "----------------",
		"----------------", X"11A1",            "----------------", "----------------", "----------------",
		"----------------", "----------------", X"FFFF",            "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", "----------------",
		"----------------", X"0AB6",            "----------------", X"0AB6",            "----------------",
		X"0900",            "----------------", "----------------", "----------------", X"0AB7",
		"----------------", "----------------", X"0AB7",            "----------------", X"0900",
		"----------------", "----------------", "----------------", X"0AB8",            "----------------",
		"----------------", X"0AB8",            "----------------", X"0900",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		X"119F",            "----------------", "----------------", "----------------", X"119E",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		X"FFFF",            "----------------", "----------------", "----------------", X"FFFE",
		"----------------", "----------------", "----------------", "----------------", X"0F09",
		"----------------", X"0F09",            "----------------", X"0900",            "----------------",
		"----------------", "----------------", X"0F08",            "----------------", "----------------",
		X"0F08",            "----------------", X"0900",            "----------------", "----------------",
		"----------------", X"0F07",            "----------------", "----------------", X"0F07",
		"----------------", X"0900",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"11A0",            "----------------",
		"----------------", "----------------", X"11A1",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"FFFF",            "----------------",
		"----------------", "----------------", X"0000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"119F",            "----------------",
		"----------------", "----------------", X"119E",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"FFFF",            "----------------",
		"----------------", "----------------", X"FFFE",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"0037",            "----------------",
		"----------------", "----------------", X"004A",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"F0E7",            "----------------",
		"----------------", "----------------", X"F0ED",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"11A0",            "----------------",
		"----------------", "----------------", X"11A1",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"FFFF",            "----------------",
		"----------------", "----------------", X"0000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"119F",            "----------------",
		"----------------", "----------------", X"119E",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"FFFF",            "----------------",
		"----------------", "----------------", X"FFFE",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"0037",            "----------------",
		"----------------", "----------------", X"004A",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"F0E7",            "----------------",
		"----------------", "----------------", X"F0ED",            "----------------", "----------------",
		X"0000",            "----------------", X"0000",            "----------------", X"1000",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		X"0000",            "----------------", X"FFFF",            "----------------", X"FFFE",
		"----------------", X"FFFE",            "----------------", X"FFFF",            "----------------",
		X"0000",            "----------------", X"1000",            "----------------", "----------------",
		X"1000",            "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------", "----------------", -- SRBC bubbles (x2)
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------", "----------------", -- SBRC bubbles (x2)
		"----------------", "----------------", "----------------", "----------------", "----------------", X"1000",            "----------------", -- SBRC bubbles (x2)
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"0900",            "----------------", "----------------", "----------------", "----------------", -- SBRS bubbles (x2)
		"----------------", "----------------", "----------------", "----------------", "----------------", X"0900",            "----------------", -- SBRS bubbles (x2)
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"0900",            "----------------", "----------------", "----------------", -- SBRS bubbles (x2)
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", -- CPSE bubbles (x2)
		"----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",  "----------------", -- CPSE bubbles (x3)
		"----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", X"0000",            X"FFFF",
		"----------------", "----------------", X"1000",            "----------------", "----------------",
		X"FFFF",            X"0000",		    "----------------", "----------------", X"0900",
		"----------------", "----------------", "----------------", X"0000",            X"FFFF",
		"----------------", "----------------", X"1000",            "----------------", "----------------",
		X"FFFF",            X"0000",            "----------------", "----------------", X"0900",
		"----------------", "----------------",  X"0000",            X"FFFF",           "----------------",
		"----------------", X"1000",            "----------------", "----------------", X"FFFF",
		X"0000",            "----------------", "----------------", X"0900",            "----------------",
		"----------------", X"0000",            X"FFFF",            "----------------", "----------------",
		X"1000",            "----------------", "----------------", X"FFFF",            X"0000",
		"----------------", "----------------", X"0900",            "----------------", "----------------",
		"----------------", "----------------", X"0000",            X"FFFF",            "----------------",
		"----------------", X"1000",            "----------------", "----------------", X"FFFF",
		X"0000",            "----------------", "----------------", X"0900",            "----------------",
		"----------------", "----------------", "----------------", X"0000",            X"FFFF", 
		"----------------", "----------------", X"1000",            "----------------", "----------------",
		X"FFFF",            X"0000",            "----------------", "----------------", X"0900",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            X"FFFF",            "----------------", "----------------",
		X"FFFF",            X"0000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", X"0900",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"0000",            X"FFFF",            "----------------",
		"----------------", X"FFFF",            X"0000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", X"0900",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"0000",            "----------------", "----------------", X"0000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"0000",
		"----------------", "----------------", X"0000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"0000",            "----------------",
		"----------------", X"0000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"0000",            "----------------", "----------------",
		X"0000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",            
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"0000",            "----------------", "----------------", X"0000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"0000",
		"----------------", "----------------", X"0000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"0000",            "----------------",
		"----------------", X"0000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"0000",            "----------------", "----------------",
		X"0000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"0000",            "----------------", "----------------", X"0000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"0000",
		"----------------", "----------------", X"0000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"0000",            "----------------",
		"----------------", X"0000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"0000",            "----------------", "----------------",
		X"0000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"0000",            "----------------", "----------------", X"0000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"0000",            "----------------", "----------------", X"0000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		X"1000",            "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", X"1000",            "----------------", "----------------",
		X"0900",            "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		X"1000",            "----------------", "----------------", X"0900",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", X"0900",            "----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"1000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"1000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"1000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",  "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",  
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"1000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"1000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"1000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", 
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",
		"----------------", "----------------", X"0900",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------",
		X"0900",            "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"1000",            "----------------", "----------------", X"0900",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		X"1000",            "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", X"1000",            "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", X"1000",            "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", X"1000",            "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", X"1000",            "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------", "----------------", "----------------", "----------------", "----------------",
		"----------------"
	);


	signal finished : std_logic := '0';  -- end of testbench signal 
	signal ProgDB : std_logic_vector(15 downto 0);
	signal Reset : std_logic;
	signal INT0 : std_logic;
	signal INT1 : std_logic;
	signal CLK : std_logic := '0';
	signal ProgAB : std_logic_vector(15 downto 0);
	signal DataAB : std_logic_vector(15 downto 0);
	signal DataWr : std_logic;
	signal DataRd : std_logic;
	signal DataDB : std_logic_vector(7 downto 0);

begin
CLK <= not CLK after 1 us /2 when finished <= '0'; -- set up clock with frequency of 1 MHz (period = 1 us)
												   -- will terminate after reaching end of testbench 
UUT : AVR_CPU 
    port map ( 
        ProgDB => ProgDB,
        Reset => Reset,
        INT0 => INT0,
        INT1 => INT1,
        clock => CLK,
        ProgAB => ProgAB,
        DataAB => DataAB,
        DataWr => DataWr,
        DataRd => DataRd,
        DataDB => DataDB
    );
process 
begin

	-- First do a system reset on the CPU
	Reset <= '1'; 
	wait for 1 us;  

	wait until CLK = '0'; 
	Reset <= '0';



	-- BEGIN TESTING TEST VECTORS
	-- the order of operations is as follows:
	-- the testbench will now load in data to the Program Data Bus
	-- the testbench will check the Program Address Bus immediately after loading in the program data bus
	-- the testbench then waits until the rising edge of the CLK at which it ensures that DataDB is driven to 'Z'
	-- the testbench then waits until the falling edge of the clock and then (if reading) loads data in the Data Data Bus
	--  			 it also checks the Data Address Bus here for correctness
	-- the testbench then waits for 0.1 us after falling edge and then checks the Data Data Bus (if writing) as well as the 
	--               read and write signals generate by the CPU for correctness

	wait for 0.1 us; 
	-- now run through test vectors
	for i in 0 to ProgDataTest'high loop
		-- load in program data bus on falling edge of clock
		ProgDB <= ProgDataTest(i);

		-- test program address bus for correctness
		assert(std_match(ProgAB, ProgABTest(i)))
			report "Program Address Bus Incorrect"
			severity ERROR;

		wait until CLK = '1'; 
		DataDB <= (others => 'Z'); -- if we were writing data in the previous iteration, want to stop when CLK = 1

		-- now continue to the next clock cycle
		wait until CLK = '0';

		-- if reading data then input data data bus vector into DataDB 
		-- otherwise drive DataDB to 'Z' here so we can output data internally
		if DataReadTest(i) = '0' then 
			DataDB <= DataDBTestIn(i); -- when reading, input data through DataDB
		else 
			DataDB <= (others => 'Z'); -- if writing, drive DataDB to 'Z' here so can write to DataDB internally
		end if;

		-- test data address bus for correctness
		assert(std_match(DataAB, DataABTest(i)))
			report "Data Address Bus Incorrect" & " " & integer'image(i)
			severity ERROR;

		wait for 0.1 us; 
		-- test data write signal for correctness
		assert(std_match(DataWr,DataWriteTest(i)))
			report "Data Write Signal Incorrect" & " " & integer'image(i)
			severity ERROR;

		-- test data read signal for correctness
		assert(std_match(DataRd,DataReadTest(i)))
			report "Data Read Signal Incorrect"  & " " & integer'image(i)
			severity ERROR;

		-- if doing a write we want to check DataDB output for correctness
		if DataWriteTest(i) = '0' then
			assert(std_match(DataDB, DataDBTestOut(i)))
				report "Data Data Bus Output Incorrect" & " " & integer'image(i)
				severity ERROR;
		end if;

	end loop;

	finished <= '1';
	wait;

end process;


end Behavioral;